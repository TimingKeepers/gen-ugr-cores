`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LjrTJsFDTf98k/CkS8kZjZ+5P2v+ejXBNE6ytIXjwXXTR3eatC0d4SJwcG7Gmk13FPUDYtwj35pE
ltPjBB3NepY+C6FlZFmmaZABPKZZy0lr8cL2H9TpyYlHc9PCsqksCtL2sZ6PJrLfnkXrEuefsWcj
fP4iVL1ZD5S/cktmQNirsGB1+vVThh9hX6LP4GgCVmZkN5/TEnn6l9jWd5uU8sPZZSkgM7WCYqov
A9HrPBq5YYe7mqjfPYCEO8lErzeJez19eBqYGsd1rLnQS9TEX/Q4jwA3dv9C+nURglr3Q/sl+fEe
ebjMnWXZ3/76a+PLdJI4gUU4q/9aH4RTDfVUTw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
e/teBnQOOdKWoE84hr1FcGfUiv8rZ2ohbbMm551FJT0FVkF/vs3duTwdHBOkp1Gn/1lbwR7243Vc
dPI61P/Ei6cyEdBPSSnYA7lWaMxEzxsXJ4Zzk3bGA62fl5vUY0/2hCBvV6xY81skxLcXWBlZJY43
yjxT9mOGUeXUX8+ZltM=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oKIrM8m1rOp03ip+lVozOz+ot+GfBoZFPDhPvnnamnbnTCx1tPnMkjUXCedL1aUaPFoaGwZWXA+7
25epm51yPrKP0FanO0yT8vPU6t8OePqCiY18RtRrzI6FnZAwXBaobI9F2bXkoFXmChcSX+8GY8UQ
2IPuWvwgitnheQiodUg=

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5936)
`protect data_block
jFcJKwp22QHkaiZlokSnCZRYHRf10PCSew5NpAuiiizPPkfyo0ktoi/TvhHXYwx44PyCJc7SeiJ8
c8+EiluqxjDwfWn15S0XWWRrRaedlAEmEP6BjL21iSbq/Ee8bGZfBN1TuA6myWbgR52ojpACsZue
WRdV+BT39eu4EmB5bEh5V/J31b6YjJ0xgX2Ey7AdyVaPt+5Ryg0hu/C2KFQ6hwIaBDu5GUUfarZp
jHy5VpNdsJb6klfy8g1BHjDkPQQ93KNIdKz2qF0AlyXH/MbcF8zmIR5lU7BgYOL3q7vP+2uU3lpk
e5qHUS5itZ4WUKz1omJF76yhifkDtf8ie9IlDDpMwYaklipRCeUnRAwTCWBI5FTAXcXmg13KscV+
8P7ZTHzvp00xL0DOxwuuvfrEgIj9zY5+uQe1I4p/RoxaFYN5U693sJjaCCQt2PppNedo6cNz6VJX
MxZY9d9XlZFenJZNkAfVvzHNQ25L2XUkXqZ/KWVvZRnOP6ICr+jppls+7IpMuoJKh/ids/gNkeLP
QQDz8L/VqkHAHad7prrsk7qfyIxXfQRNexbrqvNDVKU7mjOuGn7qlFPb2bjp/6vxN7MP4uKmuo2K
6n4KCqSi4R4pbdomL2va9ukkdX7YFWXqpQGefJDYyzSDcokFShNoSZmlLaU/nccGR1v6DIW9liJL
FUsD9RmZ81FIJBG1ahSK7RSJt/oNlyzGfG26kVNr9U3MDRFHsplZJD1e9jHH+19k8j/P7yYYg/p7
nPhIIeQqvREyR/ZN6o0up5TSYGbG9pk1gO1+53dvrwUkLklKV6R8jmRqRwjIbNy5XuVejNI4RiEH
s6qlBZZV5tVF65HOrW0n8/Hq5tjhGCyjrsuYOiPNdFPmwYxvKtjcwlyUGaVxJdwPJtQ943eAM4Ip
cXBYaR9NgQ8XZpNPFZkzg1JqARGDTyMgY++0FEn6iHZLwu15Gc6gSP4Mg9ZO6+wASWuRWuNNOUjJ
zC/UaCkIwAUCCBAqah4gDlOa7fQxks++J5UpLv7flOTWO1a5qIjumlzYtW3QuQ+0BVxFotPwD3AG
JCFD2XZPsd1fkfilsXWJM/rW/Tu6AhhrWfFFyo0zHI2j4vbHhKl8IQT9FfH8pSpHgiK4Nz6wY99g
6+Mz2Cne28Ov29099mIqsTwtlZiNz9zLp4z4TtmI+DFMSLTwY8R4b6MZXPZzSyf/DY6c3SI3B2N9
OX6UEPBm6TktnfN2OeehlDrfyubYijtRadW1DXe6aMt2UqaWAN+O/UT2oA6L7enyI3vI6Bw9OqLA
4pmhVG9sjEe76tBYM6aNMZA7zKbM5A/L51rLwGgqmM8JifNg4BLyR3sq76Xl6mbxWeqLHyGrxfx6
KnV/bqWpfTtyAIMOMi4vP/OCAXaqYU+QQ4Wriwbg+9bm207szLTfRocrA6hY1F0BrzmnsrApu5rG
TyjbIb8H3LHDpYJPmokC/9oeP60qrKo3ho2+am86oYpJqXFL6qTyuDVGm1RXD0W6p+Nzslbq4zBn
QgjG9busrVr3dygu9SvO6MfBxvieskK14n8IWlFCbM0bRzpEA9jCHurwJQBv5tgI7a4F5IXcAajQ
PZZL3nlbAUKINg4jpeHM2eQNmtl8PTZs+3TRL+BJScsm0PWoPApErO/t6O30VH57f9SVLJ90d93B
txTLW4ee4cMdw66w3ccxjiJ1X4G1by4prbGRJaOBlWroCXauCh75O4hlyUDQ0WXRSvhgNvBRuqk9
R02yhMKnT8dm45/0YKVPi/THxlrC0PP/dsG8zPYrZzdxjTauV/R4kV6GaFVl06s9EVSCPGTfmTnp
GUVHti7AuG68DBgsU0zULSB9fLghP8zjEajNtaDUvHCASbSN2iHy0jOWWVQq0MGzCu6py50jAR8z
jVBLLXHfn1xuW1V9edVsyd0Z48wGA5iBujBCgEEmmgwIueH8Q+sUw4gZzyfwUpE2JjTKQvs0pGjW
uH1/x9zE5LnKOk7oEQAfbmBwB7uvEdstzHonCELG0tLNukx/SFNpxbbfX0lFtzRKZwZbHOY3utnW
Q3IPR1B8HaHk+FOs52mD4VtBuCO5yx0VW/uuIgx7YOgO6wtkNZ+ZLskd6evrz5rSZdF0fwKBrW6Q
PIpPTf7ZOLRk0ps0/eoKwT4fFpriSQcJm7VkEHsFJ/pQBdmvFRrORP37khiWleVd5hOiKafdMy4o
3rdo+CqKrsm4V5kQxovC0BZWcQYmhu8QmVN006IMECKDBR+Aa8xV8xFUFXKo+SXyA0/7wPKRQ8Ih
tD7vu9Ohye4yIgvDIIRI1egLhF2xvzLqFacPhwb27rWmXXgN950WRl/RbjnwsIRKF/c06lSZLZXG
JldJFiL4iTyefv2ugVObPKWOx7QmI8lOmk8rr2Uw3VS2PkQLk5nyhQqiTmPNQacxi3RVSrJJNxuZ
FPrH5h7gcfaCw1uQv2yKFrPpyj0M+5siODXK3sH3dZR/9fLgDcTBt6cNqt0rpwDvSoW9Ahj73UcA
x0OWDRIR/Kgdh0Np9YdODryttcBu/4d+FYBpN6tjEBdnidQepRF/7kdPLyWcqYcY0KlZi4oVCLMf
LX1h/4z8EC2b/7t8lmxXzUtnDry1Vo/VtM4M75jvsGtQlUNiKs/ED57VtrsDHSfaBIgIr1fnJ3b8
r8SKo6uShkqItSwVBCxllrmiIH0ACdsMGiKIFwgXPUadVDFOM4l5vSypTOxBi7ElXjaFeL8qzeSN
LqxSLB4O4SmBqpipIwu0nD9V+VO4te6b+ChOTamZ/KFWAH7mubwsVtFUDxefpg3vXA7dURxND2Vl
TgE2XFyKZ9uFYuEuAAEYQrfYvB0zmtdQScHGh33+cPI7GMlm2M2ceSpweAdF8ZV3dn8wFHNGFI4s
s/ZuhN5aWzM9d8Oc+fe9xP+0T59mVhGMXnaCu/FoK8RBvobOOUtPfXMtdQ6Et+emt1y7uQwHqdcs
3rPJA5aNqN5vIcvkv3UFPsXT7faKuK226T8BtIr+cETX8paXQhKxrgCOP8o/kh8ypk8FOvUfv4LD
G9HFQyvooa0niswoR1DkSrPYydrB8rdytmzbFbFlbnIc2AV1QNam1hWerZNOr+D1LzosapNjtkV1
+I7RIvA1pkl1Bmq/Cmab7ZaCWpabjgiUebUXFL3sm17wx8ijA4zYWp8L5B8pf2DZqpvWqVn5YG4A
ojB8oGHZfMfsPtpk4+9h/6lsv+StVLky+fqIi4rDURurLdkbIH2eij6uYiTx//kMvSXS0QQpi/2y
K8JEQ5F/l+2O4KycaCAhZyM7Sx7ckiMQwVTOsi2C3wPHLNtr28evZwGJ8yuGZJlxXjuO97At8c5I
JJ+3/tquicOv4vOiRezLdjnhUBlneYg4EnwAOwlmhX71p8ne23Zctc4jRXxOAOLW+UM7Hnk61s2h
QN4CaVxwktHWAT0ujw4z1bRIRs+QK/64Rho6EEvvYXbI2qFIQdifcMus5OsWEy0+38BRpufvrzLx
c9VeaLvczUn8I4L+6iMhNGijVzQcAM4pjuLwzckNft/pgkT+Y+PBz4GDT16TA+IqjJAgp/IgtDGi
dqFvvGHihke020+c5BxkNqueLwui2xdqUZ1Z4ScFfqrvGDdAVPISWLLCW/ymxzEOnM8BNWIGMYnr
aITijXWlouKCt33q+0vqGjAfODS/cc3hYqXVZtwyUO6vBNbe8Wzh8H6oKKHQ4m7fqebA7fHjABfb
UzS6QyIw8zjsRXnjCpZKf8Ox8ssGC8nSmsAFZOBIV7StPouUBdLMd+7mmIkTY87b6tUu/4LY7n7a
I8+NOoObj0ZvYuAZh8Xxu4gIAPZA2uKLxdzcwgcAgBKTJZY/R3Wis4T33IbP5vXC0WrvqqE5IaSb
HqEFzb7RzRogypntqCAtR9GZC1alzK0BvIa8co0ByGWcaqeh+xy4R4ENyuPnG0676X3FjOVO0Qov
adUMW3AjGHMl4mCC4qbuY2yqYup0k1pIHs964gEbwqvK755myWWBpJpvIZ7hlt3ypEPAEv3YcVwf
V1tGKpBTkbQWfEQlmQZqXEvqJXiD4phd6KannYbB4x7JcOQ6igST7W8oFDHA8BguZc3VJye+Y4kr
49TWWf+7xmNvHJjaIt+qx12iX6mIlyYM4PIwHOBN98I6FSGSwi2MmGN1Eyz1Kjsz7LxVSF74JYeo
27KqFmzzRanyct+3eFmXw5BOV7WTGtjapOcUp0U/QNpnaOyYS7NC3nojhlMEEla7J/A14C7s+EZJ
pgbZTPad1jNHmHh/eira9GCNHqtqPInzlVlCKC/MX2KZzpLrXCG8W5+3Cvx6oYrQ1SX6DCZh8Naj
y6UHSmw7qLC2WkIlNlfMRDMB4hNVhf6WkXgSfVe6T9T4FoTMEjDIw9qJj749eqqIVuOKTCXZNUns
Vt3Gy6PO9NoUnIOhsSpKATnyy+zhACC9r7OCZEzT6AckouwCQIYz+Z5n9faNqpqMnw66B3iaUb8P
aR+2GAVr1EkGbymLVI3H6zS12h52UTjtdjFbXajGfWwMGehPG8IkjaBE1zTWqjN81JJaZJx86bWF
BlwmRXcZGPWdzwz9+HnO0xEmDHe8PAxL/4Bcl+JTdqxBNaakefkGfVa70W4ZwEa743dXtDXeeszl
vYa4PtdzJELDOGP3NhBf1NEvGuc17JUhBhAr4UOcV6ODJnScYqAxZ0nmgmUP1O0gt2Y/VBDPahIB
lTAQrzQJwZHSEmiTAIhokkLw6h0hN7I78VgjSRpZV1ad9RyA0XCV1ClWJt6POAe7gOQINMrPU724
ZUwmewIFXS69/uQz6u/XlVhW8alRfJ4McA5VMz9y+Yujjz0tAkQFVDzR2LvAZbYwIwzhML70LitA
yfD8VHk0kDcS1JOayJyJeZnWG+wQpG/gxFXRAIrPhMqTnoCOwougzAOSSUFzR7efZ0LkNStqFYZ5
n2XvIXTMcbcEoP1Tg7rkxGp4t/StPG5AEZj9dFmqMneYx2tlSQByFDO0gBwSm/yuMg0meXNs7Fz2
7EaG5QPSmR4i7RPl4OfvM7soc2ck2TpqQSNdngBVbXpcGMTgDN04Bq6f+CsILGFP0xPyzC+BEMo9
70+7Oal0L0Ot7xtSfvLdVK3SqazykdYd/JhSXJWN1Jv2BlgpjmMOGtydfq3O9cRvVOwGL5eL7XaO
8jpM66ydx/0LIrGDH6nco0i4XQHCJDZge2xXcXAIQ430V1NzZ+/iHtPlc4mibFkZIpdvGEv1Rw48
P+s1rIESX2zsyknMMdz3OH9PUKg/vikmlyKFOHM1gkkgvmlQov1yv0kZCi/U5riybsGyM6ANDJiO
AcwtNo3jp1wjtyVvIbKSgCJFTM1dQPLxGGtbBLFb/oml6dbKKQ58hYjBnRLGuQDzcBAoSYQMtUSU
ncBcKnL9lNui+X0PNEUT/JiheZGPgOAYE4F+/LQ5g3PlYXcmrMBndsqK68kHH0GmD9y6H01iWV+R
9FvAjHmptH7G72a6U6Yqd01IkOZ8X9Z2rKd6hETYlmLBaIXDUdWJLn+qTUBk4QAMxT6OM8o1Lgx2
r0bkS5hOMlzdAyQ5Sf91LzwWNwTRYEmT9XYOAbfc+dp59fU0T/Kx43pbV8YEbIG54KItvzOTJM0f
MoiavbBYtX1c62nFq0/1IdDWcQacCddDKENOwTAXoPSHgIkdxsda4w9JSRDN2mQqT2TFt8HlB5iw
LR3xRp5P/YCiQC98t/rs9vEHo5iu0p4ryEXt/p0HU9gw6+jIKtakPq6n3ckohql24lUTSVwHMAh2
wR7WFngACzC8QdAQrCsLPox4LhEJD0XwxkssrCZCFFeL/8VT/RSG+RcpNvxgM1SxhTCprNCx+b3P
hbqLeanD2btBVJWkcUkVJQgyvRKoWp+dAQuN3VBCZ35kUjfCiy2Mm2NmS0x6LqCgfHDCE744GL5B
iGHBWHIP1MIO5sK96/gXkepwtbvZa/WbcMYaNMjXcvQmKyFqKIayTh4KqG3J0tUaYpexU6lXRX1O
72N3jQQUhP8VhO9wRzjkN4amNoMCxIaYMG1LwNEeD+IgyIFpflPo+buOexMqlk1yNXrB+Zq6am7C
yqb37L7UdV35GOJza6cPYsxsYRGu+j8mMurutYAt59fVvcQKtXbfrJGpNGzS4rCmLZm12NOGWogr
8Fl3Y2WThUrDo2UGBBzbPRvqMvr9P2MbzXl5D+v5iAIcpRBcnPbGh3QKwuDExB3qcCKWQZRrS31E
IKbFhPQ+fp0MHXdqvqxAOXoresfk0QFlgOg2HiDRW5UTf7A3GkPmpE8gIwOlz82A6i1WYiyTKyCp
0u38PIQdwgvMjT0ovT7KLTYnphtRiAgJGT9dUUW99WJtswLn0rzI1afC5Leg1ut/lJNiqhzRC3d3
S5Rb1xnTRpZ8smPMxd3H624c18Gr3SNNQG+wN7XojxbRv/7Yzir9ylD/2YK0ZVJTCIXCCi2Cm9F7
GNArN7Ad8Q4ZkbwbfsXe7PxTfVWe4u//quoEDfyduOyLRDtr+PwmzSk5tNZFQ5g4Soekfn5p3BM+
a+vmEgFJupmWX7+LNnTTfs8UMq6Q1bBWNsrNMw891SzKCR9UtMChEB5TBgNreuiitfNQiIoifnuZ
RhIDdNF1HglBDp/MRcW+3HANvPJ/ZVKOehx1SL1Lkbp3yxCRZ4G7NfEmx2mMdj4Tw8MViXj9kO+P
hIead8jdJrgdSqUGwN4kxI01V0fpZZrTsnUuPASgPdPkad2Gx7Z/1LECDxCV+RMAgg7bwOVuQrL0
UXeyBThCkolAjDkv06nnZpxKubltYic9aNYB/CqwjxFc+tzIxasSdBbFnNteVQ/Y9+sIQAxbKeOQ
EtqBWcAiPeF8JmvB6+wfkQ8jqxrHX7FFA2OMj29dgy3kz3NMkMhvgnurk8WhIZd6l1liUmBqAl9F
pCXZUotfkKAWIWzYFVyA2IerTF3BJ5mN1kN6oK77wJCjWwkHcrbC3sEprocW/JfYVdM4zmixP4sb
zSyPdF9/qZqE/gZ6kxLkBSpz0PpkyyDRm5OnJD8SZ2S3A27WclUB5GkYW3w+5EIBuegr2ptEvpuY
9yYkH5imbqznHBFGHV/sA8jduYYnFR2XwBHihEHgPBcNT+wgNd59onImZyOwtM16TSd4FCiuLugc
XurjLdI61imUqBdcwDszSbLtG/OeahbuJ9MwwXGlGjK1dsZ0yT/0RLfI34jzoMcEfjvljDFQchZL
Ew0TIw42kZZRdN5xU73xKsrVIrdGsLkR9w21hjvqHYNUYu8VPV6xhjfyx1t3FWFq7LnG7NJ3qVUz
DnbWuKNEpsHfrNdP2sZYlHp835d8GqhADd9KrMREXcDbxqBwjdqOxPt/KZeQ+XrsOEGtaTirZ+GH
P9hQaqchrLgGJiZRGaWrCiD9Th1tgfKuo6dFYPj7pdg/O6duTrlSsyJMO4ExpMyYhyxJavplJuMf
Lm1+zKSN0Bs6pg+TE2GU4gLOU7jn+qPaRv+dhd4JKmQMV5TgmYVNkHgPSboGy6BoqivD6BGhncOj
K8KPF35qicMvFI5ol4V7/AlY1E9yHLm47Dvdw1ywm3qc09g3Eh0XSVjOxaFYU7oZ1wzYC1QV5XCp
E9ROrkpAbgvGPfHusBr/aHQ/wXhIlVtl+VcsUMJWU4WaBhzf/2eK+8guF+/TZu71x10pAYYP52Uf
xw3cG+jgmSg7Ahr8JV3H3LJxDhjAkqGFrgBnN4j46W7yu9IeURTMxFe7XpV0/KOqPcqOLSyap5G+
lkI2BOzsUCuhgEPm+4hqhHxK/FY1j7f0Cww2SrDNbvaEryLoJUDwoJN+jpRdEu+CpkDPqs1gzJ1s
60tApEUX4ARJ0klLVtX7+YfpB4lsUtcpwTdbiWidaXRZsYZZLZMUyre46vcfFza+f7c3PB+W8GbH
Y9zywXIC+E4=
`protect end_protected
