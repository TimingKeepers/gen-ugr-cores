`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L7z8De0MRldYJ4ROzPP/eLdhmO/1EA/Zrns7BH0HS4b5K4kE+siyCffRudASvIdloR/vNwAEeEPG
g3BW9pH/+fohXjypTfy2N9K75z5m7cwV5T6VSvaib1/z1JkU9ucgMLr0tEojEZ52IP+qeljt8EKO
IOFt3uqx7ki9ltCt+BOKWydXC4HleGrDhCyRzmaavG4iBQeLnZbf6weDQh1C7kdH5pGMhahyvYHJ
tvUGv+L9H3CXWa5O1LLSDXdO9RrNr/mRqkFGj5gBcutJB3Qa8aVN5HoDR0jULFc19vgjcm8wRjMY
3lcyvdWtZYC/p6Vq7qQxpPOm895sISd6nfPWoA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
I1P5YrAKrQ74o/i7roati+7Jd4D4Y/O01LdHJe3bATiHe7WlMRf/RROhErssmpbRVu6yBvoakz0G
CkZfgk2mqMssEbYqLauvZX7LGxYy9+SAASeqxZyeb3FMYsZkH3XNYiSDw4IWE6JTHvHb4Pjiwzl2
6TRA8EJeipKnQhuX/O0=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VS8QH18bY0CswpWJbOXaiKsCJ0njHIL3DAnYqVUb1CZoQ5Xuh7dQUVEvi1NSWNkqiUl9saZhZq4A
mXSuCiZzfTMCOSmVTdLF/gaAw2AF5pTynA9q9sZUDDoAJeTTnuUOa7YNsmfoRmFjeees2M4nsjt4
spSVJWPSRcfAWr+vumE=

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6032)
`protect data_block
7ns1sb+xYU8KJ1XArSD8LkGK1Lx5XKlkPVNbQ1muUxBFWK8vlxQYWFbQkQkKNsn8v3xa5TTjsIvS
eysCHx8SvB1xOWp7yX4dlb4aLFoAT4rfQdgn9FKcH/e56SNH5tZNAKKmOWgEc4dNbMoDaRds1f8Z
AXZrHfcCS2Kj+9sD9/9IN5vhSDb6Pcn3BAPV9DQaDbhFr6WxG4+ULkoO9hb6lm1ayi5sxCrWpgzv
3A9t7AmE8+UqI8NwC73F2R2YwUuAmq6KBPg405oDyTX5YegoNl0JpV9UjIxoTWXKXPSqnU+2J2ob
a8Cy1z9BC1Cas84NrtIyXDDy/9sUM8oPU0HVHT7rdAsa4OQV8jZI9azEc4RlTmn65lSqO2mSiZao
574CavpmIHn5P4E88/a1nP025guBMHNfTJ7br9Lt45oeWJMCEcUgE3ifGhfCx0q1K4ef72gKFyHV
546j1lpc68HXY4ngje/I3PUE19ynljLhPPAzsTK/eq2kqWlfOekaKqzdD9jKE5jtdoFRwY9YP7Og
SsJNitEef2oqGI3u2ltXqfIVr390I7C78opS3B0xguuF1LR72phG3x81SA3pc+zmqv1ZUaY4ivmv
NT3NY8139KPnMoB3Mf9fWp2j3yDfF7MLJMO+DmGJ+2vKpXouxj8ali/1CVoYx/d81SXXtRKJGYbf
b/I62OAghOOE03iojcUwYBdsjZsDJI9zKLPQmxYvAoWw8fImdGUbnvLgKeLATn+tnTw7mUKdtEng
GtArHaLkynT+aADPcpF/85vHFqYsVSHFTL5Kwqfs0GpU0paIZr7x5twTU1Nb5krPcVPwmeV1MfQT
Rk+4t0wS5b3OUQaMxlSGKHgYKotgefKjw12odqaSfJyf8Y6w+TZRZ0rQ3o8jyH36Bl4gkd82Bb7q
JXN9laPACoAr09PFvt8lv+Tcrkv8LyB6lA3e/l3+u10ja90+Jls3O5IkkHaND6BIMrJifvv0u8ZI
DA7s/+L6qEQg9hPWipvvaSv646wKQn+062eDnhTQiN6akWec/Dn4O7ASGE1RLwrsRY+4SZlf5aZv
NPrSqZHpwKWX1IGMGMxhobm5Bb+tbiTUy+DNItL9NxDYPiQqypGmKS5EUZHWVg/N6Aaq5MJDUzPu
EPo0abalvs0nFJY6PLSvEX+QpKNCM35TajJVZsoWJ84Lr8i1sW+qjQ2aav6h6IPkNCWlCPnc2YDp
JEVY/zom3Yf2KVymaO0MnaF7fDzXPY0D6RuiY2b7AwFr+6BeatKMgVfX18KftIpFguo2ZFVgFsQC
YADsNGM0z11SGkeZxV6FgeDV5cvLePBTlpWdcAUQjWoQf7GI2JPyi8xQW9IlF8ihL0ZCvvVYod3D
OQb5Kv8DBecX5TREHPVqNAG1uSTQIqXiZy46Sv2+LG2lGU/04q+EaG3i2oYX0TFZYARinWReNfV+
OWmAjHC7JipEPflZFScDzV0Zh4mo0y9MPw2JZ6FKYPtbqomllOiAK/3wD7pYZ8hdjHfIxwUxZh4J
jWZyCWa/9qOYKFC2ROFJP92s6e4heSzMCEHZCPmJSdVKIRlncSlHNrEblZ1It5413HIrRWDr1bBb
kBbpgI3obV/6GP8NGARgdC41qHkLw9kkeKHB+Uekemg7qyiVL/WwMnVXPEiQxSPA6qt+jR8YJy1d
zXUO8AY5/6dUK5J0CgdDubCzG9kten0iCA4yNai/JtsjtIlAMKgCnCX1K0D1xuR/XP5Ayf3XsQJL
St3oxabPL59Stu57R02A+cy4I0XOn3cYKfZGip0rEpXqFemSUDes51mvQQnv6Gp2WcNH6aLpGwbn
m2vNG1ZcKHaIe7H93g33I1qIOTSg1eLmonhwEXBri0EwpvXkxp58b0hCilQFbqNyhOfmC3oLyG5B
jD/iCRrDkRbA3/7T/Dd8cgyU+quzVF8zfbf2JEey3Ui/w8HFJ/VqWSBiICKEjAFJsHVuGMyJyCf0
uv0BomCgbYT+osFWjXIKrSCCqLfMk7BzKoy2LYviw9yRlN8lJT9eMLHEKzmNsvjG7FmMNOzdtluc
tV377ZfXmQdKcWjuzjosYFHPuZk/w+JHWp6Wt/lBfkQ7z+k5m8V6FePo7rwkiRZkikLQJS9IN/Xz
62Av7I4LakOFU2CEf3nF9o2FxxkaMz0NneRP/wl7muyax3HqKVSfumeM9U6oaHfOLxngUDh1Ns2f
TboBfyV1OCaR2NC3l8HpDQK18lzvJkoF4QJUh5U/WTq2ke6aDxIeuSIuNx50rCgB9DyepWxMLNIM
nIdBMIwRERecMadz+E8+uXXYs9eCst3iXj3nN8BBfDawsahdOMWxc662hwETLwgxqC+3irxi2NiU
Vd6HA9FWzvDzsueoD8hiuY1qkXXN9KXm+h+FMYnFWpV7ax9+G/i7EovJueBT0FzXyvAcnhF13Rkv
RJFTEIw05S1o8EbNV3RTW1dqsa9bU6Lhk1XbX0hwFnLhJdMG/xz0+g5JuNkWv+KMLRyVroIfMBjR
P2XMy/pjStC+R8KbndYFmAftamPfqADxfmYzhg12D5qaLC9nndy3whOr795p3DrD+2knDoqhWl1d
J9i5Q49IDaDAHpfAQEcok+1Pr3LvcPZ0MbKo57//EELmmDxabBXtFkyFTR2Z4n0jjm8lJrV8riXZ
LFTRMLwJWQlboq2GnhOP6J+pY1rqF7c3vrl+pt4s3q3/gTjznhv0GSDVjuyY/hpsXqxNYTVDvigC
N8ko6fqTN4+PnOY/01UsubHBBkQJVzwBGpCZQVSzbYdE5R2zMN2c+h2MQgTp1J6otG2qW3fEX8pt
Cs88ma+NKfre8zP3MEAlZY1Ob3QCAv02ZLSZpHWmnImHPoItWjqTqsQMccFysptcl51KBhJBLtsy
ntunYTqZlb3ETErOoZoS7op4y1Dwkfvb7RdQMYgEuuay5coNLVBuhlYgWhh9IDykg5Iqcj0W5rZ9
wMlm49BKeEJh/h9s0hMRyu+CcQrOjYqvOEAAW8DsH3ZkatAJRf6rxg5KxqkhLchYs7hSvctZQhoZ
Lxq1zHwdu/uNrI64DB+gDn6wQ7oGjz+LPF63snrYy0lNBD0WrNwkbLljA+ARHav5Kn3II5vFkLqG
c4qevhmc19JDFhEAcisKgj54SbmExrOIDXBmV7/vtraAQvm29t2Ac71q3MDUPoVOM8/cUBKHGRKU
4ucMnMdDdrhzpj527qgrE5Ornk8g+dWI5UTMFezkq01s4kfeiVDY2pxkJ1eZXzCra5mCDbDSv3et
LRl4y6TWiSMF3b3tj2aEWdhmL+7lJbCfp8ni3dIVmk7p5zuNk2GnnMhEwD4fU7k0b3FxhUB4Ob5N
CaKuANNNLSDbcCgSUESFVs4PZp/SkrdNWzV+Y+L2N9WzjNTGl3L0jPpLdr+TOfu+wH5Y7zia+dzf
RsdbpMVDVJbCWiGX4lsVirMZmzv6ftq0hlZ8XgCeJ+8WOyZA6B4GwAh7OD3izAGH9ZSHAzts663b
dEArXCgN4sW7QZMd7e3lFZeVbHPQunEyx1U9UiK2+JiXaityx2hYq2l4+JoXqx5CtGBmFWl7T8ik
iFTznLC35FQk2YDLEjGCwRDIkUOqhLqUacnW7aw4xV4PXILbcwk/pletsiOsqNJhJBIhC3uWQZNl
pUu1fbc1rwpUGew6H2Bk08bDJzzMZxN2LF/WVrTEJMQxGSSc3v5gSthBMNTVMo3//A0Y20W+UOfW
UVO4psBGGBqdQE0CuQZM3HfAp1awTTw1+rYsHbM17tLERYVm5mvW4B0nBjRWVbJksVZfZiRAc9i5
SSzF7TLvU7znXeGpqyfkUZjQO97d/YKYhB5eOP0VfiUhN50a64lF/iYMJtwu0p7YhK2cDRA5AShB
ksdQ4rKXeLBn+wURizkLuNw/IXsq+T7SB17pNCuy81isZvxsI+cJHDvo5fckL2nvklaPw19n/PAr
e+v+wZN5lg8BGSMRS9J5qYmj0bt3U3Sw7p4qvONqW8D/iaoSIO1okFkFsFemtxx/UTlbfsLdIflA
7JQySDQNcdJAxzkK8XP5X7pC72bGhZfcbPgTXw3kFmMRvVRRuf+cLsbJK84jcc0O62iaQD8dZYGM
ebCesff35igW++UdCLD8pgHJeDWMjoHeMueFWG8tCb/edciMTP8Ejtf/ToJYz+B+ekacz4TSSZSm
umyXqgn9+S7QU4BBFELUUl5D1zXNfCkJpEXEzVMC4jCp8CE4a8lQIW+mZQ479c9qzy+2gEuTIPdV
g9+lB2xIA+nYoQSlTj2neaZC9CylFM9a/QDzt88Uyk9pahDJq2E7vZuP2tgPZ3a2GwhWPoD7+MzJ
rCiA5bTeXnlBuV5G9uk/QWM0b+cBLLCzRATKPIriX21UxZWUhZcjlWhkjR1SMjixQ39xIvLuUk3J
wGwr2rE97EP4mtno6pDcgaB/PGl9RFmoFD08AoySSUlGBoxJO+9TeZJFtvjv3VxVrC4NgumQ2hK8
Ld+FS+5BgHfXtKWwXhgLUQAMNIQzULtb8s9IvloW6gJWrz01p6gLIU+tJWhZyxhgU6Ytady5N+Mz
qDih6NDBCsnLBOE80KpPLN687A6NTxGPwGjx09mg/nNNA4fXHORt/2z7Bi+j1r0NQGyCuTrZ8BB1
H8MB7/nO4H5iAey4it0vnydSx00FmXuOHtC6NNqSUXYARN/Lk8RlO8CgU+DtZZNUbZcvAwOHyniZ
FH2wASTYE+KVf1LemnyY0VUwg/00FFsvtHzC8ZYKl0qs4MAxKjDuxLlQLPOgNG/1xky596maoXob
QD2k+kOg2Y8eQrEqyzuIJtEuaLpxyCp+sHWFtMj9+Wwgen/jEGuNWXc5PQ0iqNTkmZVYuLddopNq
lQpA7u+JGssLYo6JjgVkjfw8DCEhdU0SIe4LTTPNU7ltpjG9wCrLsaLAKRSgoGSKQmvY2b17RVyX
EP6bXyulakxMk2eA9Z8gaV/kdzaOzSa5ZXOVT2/9WI3wPnfgzBgpl/CO+ou1xiDS4EkzKVSrQI5B
ortQInm7IHmBSRmiNuRfI/kGP7zyZZ43VKxbYaaeh62T10sXxgrF0ziSCJlrXOZjmdliLYaC8ITg
KzilO1BBi9WodBs8PB5/ZrwkzuJW1BLvguASSFHDVBvE4eOjmBiWJ0OUb89oMSCKOGRx7qKR5Mg5
3rOt2KI2N9q76WJq1Kf6OPj2mVr5i87jdToFkaar/VI6IOGhXBbVNh36y5MgFxzDU0EIMrW8nFlb
bHWW9AYsqMOicSEsoLq87nX/NX4yvGajZhLi7Kf5IgFcM5xeYNyVHZpbCOZ7qcPrh9SZifQU4US2
jr5RuzRTIUIE1bxaDq9nxFZ1ipa0ETk4RfBK2ALv5wJVdw+NxDHlWWe/9Zedb3ozrHWhtGSIri2N
7pJ4l3o2fgH4KW5ZQQ7ilsO6C6cAOXjNK/5AV1ouH8o9YETTEYa6r//Cvs0oUeCMeF1gGrqZcxqy
ZIFkWCIp1SAdY+CUpGkEA/8wpA6LaE8NjuX35U9xF4IJvyoRgoAZBnpm3b1DAot8JQzEy12/7/vT
Pd3b9+HasseVQHlLFsLPZZNZ/TO16GCkaYbT5wNk/IF63UOFFmUEUc08UHjYWsYox8wYWJk7naEg
ynKYYK1rwqEVrk8IhJ6aQDiVNbkZ4u4IkLYr+2dCLeO8O0Oi9FvGnSXNgYByW2lAZC41th39JJmo
Nkp6nqUFNKtlxmbOB+L+maY/fVZjlWnwGVj2s2csBzPA2YSSog0j/VZbXu74BulaqJNe4jUjGotr
8APPLdatCP8zfJHNIFXEzErHeUQ6uDM8lBD8WVdZSC5D/TcXLffAndZ67/k7ilChZPH07CB0mihK
fkxni9nV7oqWUfy4FRkXYypy1YgUaXIstjwz2NOIzlEm9LjxQCUxdlkvjpoS2bnaNzDNGXO3KWlI
+8qBtRRDTgzkv7Y7Rs3TLf1k8u+6ECw40ZJWz9SyuovfdPy+SuwlV8OP3vu8OqiKs2t91qaFPcv6
BTTaHu8fOkk+jWU3SQjZl8D8ytH6BHGrI5R+A7NyCK1WZf1cwFjqHx8c+BFXQe76zu2wRlWeTRaq
7OTrFfhAIfH03OKlkTcFMdjo/YiqM3saz6zEfyCRNp76sdTh6EL0uYyXYg/j2b2Y2wFNB/QeGdPL
N1mOaLN0/VOEEFXs8S7w/Gmv904hmduDFnRVFvgW7ZdIAlzBHicDiDBpr5PdRVi392JSxg1B2mvj
VuCm0CDNnpe2vG2hn+ipirido+a0wZai4uwgTWktqhH4Wgr62hzTIQwlW/hitYqxwit6xytgA7m5
07QvPOv7/rruM+OXGsIeIbYHAY4eKj4HfUBTT5TBasfHP5NG7kOyKOJ1wWeNRMAzczzCSpH3n3Si
qS3avO+a79WiabaPKsujDnnE32GkMl0BAkmAc8XUG9zNpmKo4+/U+uKxgZ/vEz6dWIkHI33D7ijv
+RZQYQx+g/AloSHZjbF8y77tSEa8XzILqLUhihu9dETSYqSzDWudyDkLt8KTUTfDZzVSUuKVusEd
bKwlnW9sL4ti0x6OnHFZIujXoAC4kxoqg2F/teQvZlX6VNF76tcfSLio9VQFDQwiC1FVKLLTVq3N
apnyrsbhjhYLbfSZRHI3KFmdGAh9kyat415K/yV39yeBIDHCriFt35whkO0A1B+VxDrV7rjcjgRP
HGW/rKmb9SEoCjaB/dawVjI7MKn8raTmZNBE1HGTbf0zdhMwEqMy3th1YlnlXQQtQ9O5Bgy5uVEP
NZ2Oxz6CIl5CAOFYpby2A1eG7YoO2Ke8feUZPXVZtUhujDqkH3ltbtYFuD/j4G9cwIP49IXgZbBm
mOhSy6995PKEjFk01zaiLqSdAbEob+SmA6oUgx3q0D8/spxeJ2CSjgvGRODi8JyNUAsK6Bg6q2je
EWS4/CSEK0hOiIJo1tXyoqz0LWWyNJKPEEGK7tnAzsrUICzZdYDQB5K0OYOon/SU9HwbAwrZephk
FkEa2GENd0+OzI+J6heryHUfmIuEIe/ZXAXwp8hFcjvlNW1FGXJnAN4tl4hSYznNMM+FemfvV70W
TwqxOkI+Q8WIsqgVXIbbbfcwFqRTA2CvQr/01XVkY8xWOnFAlwxk5CI2fmwytyvBVzDYsU3SEgQK
s4yF+qAAtPGO1XJ/EwMt9qGqOx5qwmX0S4+bDKVE7RjldpNasfVkrjgD+KhzTg1NUcJQgalHEJYM
aJojrC/rdeMXh+CMCSnJ80DVwna/mV8OEoGn/oaH5eOWdwdaPUcC8piP/m4lJbnNvqF69txqGkhi
ZpDvuhvTt1OXl8RypJ8u+rkjDB48TMrg6O3xKEM1HC7VqT0VLcSqpciLEd5ex7T08xJ+mGMN67Ff
ej+CPxINqJFzoaNDlYy0ouU1i5ScGSuEn4RPcrb+jHJwwaUZ3WyYahJAInCKvt4sGeHFBZdZj9LM
3A2AFg9ecSNEssRJiT21TJluHzpkcKl06wwyM16H9TLzYABKwD9U0ynxnZgc6LACM6Qsq0IT5n6t
kJZICJdH6dXGvsv4CzA6nLpxfFDstA+Xip7ar6lLtrHm6Me+xxUZQzmZKEJfsmtXezfjHvjCBIFN
LTAy+ETjG8Ky5BLzE6xQ/MmyX97uXTqD4yJDtH7nSAON55VPXz+1ZTWmwgXzy24LfzXDuW4Uuo+J
K6cAeZCQywmWzQ99dsl85RQWQ9XyBSFKrCNQ4Gvk3iRhzRIlvqoC7Yxyf70ql4JLQJxWjIxS5lEV
SpeTcdSKRXvPrWpSwLBzRbi1oGkEhkPvy7zPwADd8DJJ5a+3NapiSNjSCHTmQ2pEndQqhyuny3kS
jUeB1kw+oA5D75FEx8TwKadnqBrEzDDwunOdhYSk/lygCGj6CR1rpDh29239aYxEZNoX/bw4gavS
rHdM0+lCMlK1hYxOXq2P/J/M6CCo1N//UfukPtygLto37JgEjWrtPclYw9kLixPlNpCm7jqVyOUq
0jo9x2EYe9Q2sxfipyMYtdQ6Rq4QUg8a+iuS/pPWfbhXKeTa1vJwELJAwkCLTuA=
`protect end_protected
