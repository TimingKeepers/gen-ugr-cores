`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
f11/XoZy2zwXcm7hiAQZysa06yRMbVpUZJxVl9YMvCbBlCiCn8ZZ1DW1OwB5msmkWwvT96HBro5r
TUD81/BAs44PnJg1Pb5gPD8eIZj3JU/+so8d0SYEhJ6ihdDjqoZwa1BilqoCJwkj+rkV3GsM+8ie
kaTxwoKMS7MbZrYcx4r0ppfd29z6pgwKUkN9tdzwvPuo7AZuJBrCFq/bw5FQ7Dxcmk6QhU/4j2kh
QuOSKOO5D/tsgJ2St1hbJPrvxwYANciFm3xTUGV+zcTQHtJ9JQ0P2I+yEWVShJSMuO1y/62eu6Kp
0RYNjh9AHTNgCsoMR0fZj+w99Dc9LsnZBx3Vvg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
V184wi+ffFrfmzFd7iU5gqVolaERJC7g4v9xPdCkzirVUY7nCIrdI76U+ijAngu6g1ytSEMdJifS
leerv0moZ4XPx0nwlvyn0IxLoWPGvrGatAztH4QRlIRvt7lZYHixxYe9NgGbGkoy2/Yc3ap1v7jC
cGCu0EbxnbitFuQ9VoU=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MGplkGTKCVkz1bnwgdY8SZjAFlTuqLPXaKkzYo31CFGEMdQFtygvOor6WVEPN4jzedbCg0SETuOB
uoCp/fJJ1Brd/zNf7eRz43uaUfGZwOX/XtXTlpPvQsbAlPgHbaWx+mmO5ZInHNy3j/dznhSAGGWz
3MRxh8iQze6rddY3A0o=

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11088)
`protect data_block
/vDoevVUnAtdyQmWdC2DC/ArbqLUll8/oWAcn6syPQd4qYyhWunuk3ubEOgP329XFM8a8S0/EbiZ
eobQ+GmKENLgsWejbiEQS1hZG73rwdv6uWZVPf0w5WJNtNslnU6vXQBcc+vYZ5CQN0L4uICOpqzQ
JkSXbZGI4u84CR/eoGvgftuRGU/wJLIeGGsBc+Q2QHrr/ufzeYGFnCCBoI0xqL7vhrZUEOsQUU56
YQNyLhqk0MORIifTMrmoizA1HKaU7TE0+4Sh/yRGZp1r2za7niUM2x0g1/D6xuk95mr8Xd6oIZGr
H6tNUBHGCmvOQn3kW3unYxZqX5HTb+hEoHUx0/+E81uojx2u1DqhG0/Dv9yuK9eATYHdNlY3VMT1
mtEsMPsqPefdewRL3/Tn4QGmDBNEPzSEPbt5Yc+qlaXqbz3TuzDI0im504aFCkxFeRp369uNlE1G
fNm1QguOPVaU1UhRIfqxJdEqzkX2eNsKwF/5YZRSIe9q9Ghz3POrgiZVXFdo8rhO42L3athmDJM1
oWOpgdZM6nT7k0cf3c/kg3Y6Ef2iUYVNpwD5CEqpdfQqBMfP12M90DRb8359U45I7vYMCE7C9sUq
3FX+KrMD+uFu+Agd9+qwN44Mk6R5N1Jof97efocW13zvzWbsl9lG10XWmE/3UgMtzi6x24EyCZj2
LhviflzLCItJ6JvW6BIdMCvGVJCSchEBQ49MjgXBIf++KT2GYoki6FhyaOMUCtEHSy0mZ3u9CaDS
q0Dh4749s7FBYhg9eZA4GrMAt0l/OXy9gFqdBl+08Np9SsCBOvS6WFh0QY2cu7lRM+Egelkb5Dh9
w/aV8IvItkGYzOq7xZYmfWz1Jiwq8TODkbreVbfpOqYQhnJETnNRhuIYSCfAV0WZqvRfs9eZiMi4
smqJ7Oa0hs0FD/ikpk0TAkovAJZy+dQY6bnjvyunPbH1lsGDFzCAXfhhb740IkjZj7xH+aZ5fQeH
7ShnWHHchPkkR2U6qyuVoHTRWWhfVg1GKk8oGoyclktDZWCcIEAV+T19NaC8HcIgKJpZ5uoSbrPY
xRnD48YIHr1uLrtGkVVaISk56YtJZDFyOweo1k4k0E9Fb8BOzxSAk31zrxSv6Z8d4YKD0Aa3Zcbm
5NlqgVipdkY1TtzCR7yVYSvp/73Dmy9eZuMnF7lW+nUP04Aa7zdHjt6VsctOipV66er6K+QgOoAu
GWMhpL3sw3r44f5qLOanA95cWW2iFMmWNYu3Dfl4cX1Yn9ECwxhj5HAHSaBibnggGIplLK94zn/o
qz+unt9JOmmoKXhhL3iqkO/SMe0+qHN0ik/v+NgnY0emu9mRhCu2i2puEzBN1NcaB65AwvRIS4+j
Ug3z3mvqMvd/L7EJ3bii5GQFVGph6+KKMIZOrDIh4OOxx6GcwiqdnT+MYypQoBd7eHSZeGWLDqNs
agIixnEmWTVMRFr/4EzrIdQXCtOfFf7Q2jwnzaipBCvOz+Yyw1NM9+taWRnouq56mgeBsrqkHSXo
T4aoMVsvvrv9rnX17FXZm2+/euyoYPFuhFIzeaU7aj2pRvllMg2oVAmiSj39g8cLT0CYXFbt3inW
7LIWUFius9+KPk4RHhEfk7KIDBng0R/QP5UOY0qDC1TftVjcnXXGVT8ap8qccx4ARxMdZaF0fIqu
gMRKly1Mczjh94Hi0050PBNtGwZD4M+ajNR4n0KPVezDriZf4eBZmUhhQUxhWSnFTNrBiB727ZEj
LW49TwPPGjq8Ca6ZU/GKmCz7cWrHPRguYSyEKXJ5pBjBA6o0TiYmGwcrc2u4OQG8m3BE2GjrmwNu
UlWzBIQ5PwmkXa/MjoYqGyebdnHXhmcQbuHSEuM97um1jefchF7ktrffCMPV/D9wK12bk0fAgH8w
OnkHyx45vRfkVdx/X3mlkpC/I5S19zp7hR9mIqDK4gWHy+FvWY9LqlKSro0DSLbO7gVAF6Tx5xCD
dxapLqcoueUacaOPTIr6yn+ndAC5agg8h6rRGC8/fV9Sxl/f9c5gb+vruhjsMiXuIJsB+bS1p973
KroVU815imT7ncfak7wH7sbIc7XFuA3Q5fZ1U+enpqZSZF+IjXyPz4Rh7ns+uUHeXzXlEUrOP2Mt
xcl/K+BdQx2lSI5Ia+DAk8aqq8F6rwA3Cme383ckyj3ljR4kZSUaxi7+6fS6e+sB87Ut7ocTksbz
sYB72d0JZ0iTZET7nZfVaatSV+mRZ8m0+c7GzRyeGWn5xcSuY1oYnKZWaZVqOfw/1j4fojiQ8uD0
XFGqH7ld9zEQkiWlwC9qMdC0obhehKjtICWHpBv1ZeNbfB+YZmvZQ+L37/q5rwmEHBRR5wdUTDg0
mCo83qjSiMHSWfUDMu9Cc0TNJke6WgiR0C63aa6yYyJF39ne5QCuvro920+SB0/L4lc5KyT5XVm8
OnZq8JO42pjDgzJqNXs7vAFN07EFw+FUfLW++jChRD6yJnEXH97tXYMWBOCKI945zlSk8tszXEzi
spfjEpGyMJGKppdQ+uJAnC0sCLljehWS8BC05/Yyzn2RH3PoolwTwmEr2DJtjdFfDfeNz3nmQrBL
70Ajg/2oZ/Ikm5KVezuXHMviFekGow94YoSGaG3cMeWGkWr7ndxhq+CW5sFx1PMvKnwh4+gA6+4L
uVNKUw7GHLSNt0YUoBHOQdkn4eGEFu1oM/cLyUTTTadWB5huNgIkv7BAjDnzHMP1F4l9XsqWi4W1
l3XqMKOP++FU4iGdjHDpM87bCgwV+ljuyKynoZ4a33G4R53pVR6wNuLSyJmv3etyQQ6W0kfE1Dou
PU/ePkP9XZg/L4jvKLAoOa1pjsLl20X1/ZQMNXHW6ZAN9uT01YQl1BlA7F1LOSbdw5EdMRZWEUbZ
heZ0B4c5rz+njpVs9RiW3z3H7PhPs0MZ6C5Zl0OnM78KedS7UthLnXHfQwaCoUo7S4n7jsb9tDuH
gurZaMGVKlLHqSM8yvyaT/3M9kGnPkHs2AvC8eB5av9lKHFVAKHkEQfj+jDRpULCiq0dY052eslx
XeFWziol2YLpQnOQWXqtX3J7dk9LzpPwnM8DeL3WCOghdwYU8XkxSfLXDyt6kP+cC/feIi8qytBy
Ye8PQpx9OQCe1VFgUO71cBvVhFYfByZFw7LNk87vEHk0K/Vgd49T3g5VYK8c/qKtyNUbDxaimrB7
pOWSHNR58UhVZS6Q97VxmEeKXfmaQI1If0ltCywXrhfIxQDOV1HWvKIYZBoItBhvZEiQ3OulATRS
HC/33FmBIjqVjxwe6BBm+q1Jd3C+lm9ezXH/+/B3d0PXE2Aq4f+wtH6dVN8e5ZGH3DfqKyU8DEUr
jXQzYtLatgxu9d72eI7P5MMBTnJ+E6Z9y7AyPFmDUA/Nzg6Moy9X2GNy68EbvY1dv+6x3YhmnG8Z
mIvpxmmQghCzoc3WFpQhpZf87d24R+10ci7vjQssO3O/k/2zTjcKmILSJNrnPQKAIaiIBBme4PtY
A7/t8UVTSKB3wQJJlmS9k1cdHqV725mHNXU60BNnMMPYIJZ4q+xygTLGgwL3VAuoD6njqE3q2x0X
7Kit/8Tzo6HlHDqwOwiVMtLJhgH5Co8LJkL4gbAmTKEThqRVn4wCJLn1OqI+HpqYJMQH83eZBHTM
Ub5oiyHyOhWBcsplDBIlaZdCdRRArdVSUgonpslefJnSe6qoqFI4PFayrU9zFPuHt3+vmdy9FCKq
TkCZKJ5kUlnFrC4PhjdaJMcWoIOKpeWX+yvlWBlbSpSfM/mSVdQLZ+mSDAGoAuzW4kJNvhQ8HJmF
OCwTQYqVvza1dNmt1df3UhdAmukHP8BKOM30N1eNk88pdTLeGoZAWm1+yWSHst9FpAZ8a+3vJ+hz
nzbfwJdjNXWMQXM/Q/6JStf5jdAElEnBOVvmGkQbmllxUf8tet+46N0Wm5LsZ3Xqy/dHxc5SPAe5
Hzsdm2mxMC3/t2w3mO4wjcmZWe5xb83ycMFPz4g7Eax3+vgsg/RJVcyEo+Et0LEvaLQzCGDvw10Z
jtvA0+T1YLsX1lJBI84nWOqA8UOPqwfopqmCqeC7uUwlIwEGIpX8wOa4tpODxLvsuoaMrvbGauo3
rzheHAI9F6muEML9ZBwGl9JCTmZokf33bb8bSqB6aj84+1w0tYUxrOVRBzkArluUInkAyBheoRKB
0fgvM8qorR0iyD4Q0ipYC1hv4RN7NIAZAc7eSZcA01Cxl1lEfxu6XedSx/SbtBVbGPglUGkD5kBP
wh2zHfF1WcMS9d2ReU6rD0xsKHeCKKpeyYmlSpgTOVSGTeDeBe1JXbHgl+ddgmScnV7VbP5WrAzt
D/UqomMwUvIEsnBmbicN5fKv3XBqMqx+WrszkjgX83WMBpksGCFoWgHpyONRpzolJvpNgAeYSdMg
9uKHtSpQaAql6SdyzWBQef/KmMIKSZ/Kjz1aZ7Y/X3TepMzpCqKre67XR/a8xdWR3Xd71srufhYi
NIjIWN9z0+ecU9mhJmHe1w/IjC2Idewuf4YKgksSCQc0cufpBFzw31fD+Fv9JfO6JeYHCnYS0PDx
vvLvq5mFLqMVSgQ8sYKCIewBaeOTO1QKOzeZYedqx2JXgFhnzfQ5iSQM8s7pjHVl7zCGANi7j3yj
iUoODACV6PgvwerfgfM8fEkmGjbt5C+mxr2QrmivMofWAamPCwIFhIiQe0Y8ef9KP77Mj4YZn72m
eENZx0xXYh0lboCT7+G8HU1ArWpdwffrBHX/69eB1zcLYMoQdCysKXRoYXX9H7eotzWYPOkmL0s3
lkii0gZN5wzSVFH/lt6qAkDJuFNWE1a49ZhK60OO4LK/SXUYqLx3vbG7Flp+EpzmUG856NfVjYeR
7M+C20yWsgXv4Ac6NHUh/TnPQBHRCTyWgb881qNbqfRDhsYE8ubJrqm66qZhQ7dMuW/Al0l3VRbd
DsDgkuJ7E1oQxpgb/Ze619tVr87LsvgePbr7+o3ffqI98J5Jv4iXye7j+//hMgLUymHhJBwR89FG
3eAceUrG8JZDPkoKm7emfK44Yn6zneG3o8ZT083BHxkHtX+LNgi7l4dru7Az7h5N7fgadwijG9yP
wpq83Ty14QDQ7SJmxbmWRTCo5uUdBa3Qpd0Nk/44EjJyMD/EQNxxLWvv4gHY2UXnYgR+TYeBUWF+
FIv+Ud6gX0wZYFgJ8twBuws6+CrHil7lDvS1Oj9eWwikf+NUFr9UqHsxHoN7Dy1sV1lZyB57+XO4
18daipP6kd5bnoyDBe80+VWl82cptOfPlyJYpHUg+4HcKzLqON74Gg/dHyptxDkI6IGKzEHVWoA0
lr+CX03oXY4L9XBwJeHcF+sJEBL7qnC+d21SS6CC5bvWo4A7776GAeqha2/NlZEY+Unx+NrhMg6Q
P4Grtb7O7K0FCLJ+40IhahjpDHIWLnQNSNmPpY++m4BQ38Z1oO950SVm8pM/es24trJW6q20hEtx
/yMKJm8Eapq924kMCKcLRni2VHFZ2V96Urj+2ALFNgJOaTaI/2fHZkjzYZh48/K1DxcOn5MPbpni
Jdyj5gdccHS0fi0jAK7NamSjiqOejIGVzYZqdCiWL8TNKZgwo1W7yqKWrCullQ0XfZteDe/DZjCL
L7YzFmdD9zx021XAtJeV2X1Zx2EQ3RVKWM9J3IoBBc6DXDbVJsRjoPRNxJ9WBTgkBZ30m1T2tNEU
SwP4uCMsFnSgFu8ZQuSzMySoNJyPZPPOlvvSCz44SBD85khT+ehM8WFg2vm9ezl/UL+hIw4U7N3L
7LvBpb8PAPFEfrCvoSY/JsX4uHxI/diEGhRz9MvYSAwGrr1ENpkEtXxfLen+s+HF2MWMMLrnov3D
qql/5ufffDE9mtAXpJ3SQHALsJ4cuZvmpQvSq1AgZbgR7bRBwM90xda0gL+VTG3RASAhXwWDEvS6
y1IeMWR6EzcZl0+AybVmSGtDUfUJJBd6KY9RmyEWi03jQU0oeHqcA70+RRaZZ8DjuXx6jpzSdMMk
05b6JbY913QsGCMlTLttyi95TxHCL0aCbz0vNFwG1BxjzQYUWzQRRhdt1MKtnXzqXAn922xHcEdT
01yeoO6sAD0DTS+stlnB0RRvz9ntU9DeCe6MZOub5RCVeCPYMAQkkmmW7PCYJvYP5BvrXcL+hVSe
54kLueUBlTQbUa2kShtIaiV/XJDpfXJ8SwTpXBjfiWDDj74irjGpeZuQgnZVNG9Lm8XL2Hot1ixU
+jFzsgoG1Cuf2yCfKxkUWbqQGX74TpSpBPpQW/TCEtvf5+JT0VFEt2t+4TvfIovMcuO/5568XuDW
KsudtXqwzYFLcHxbnlqMmt+zpLeEl9KuLTILxpg/nlbGhd/g/MKwIey14J3P2/NmYB64eu/GbVyt
QdApBQN2zpjiT6CeIwTDuU8ncLYKsyvOGnPu7M4TLFjp46FuBUPf+Aa3u9Ag53ZRBwbDXXwVy+Q8
EJWbFWJAFuSrmau2PbneqQIYC6LAoNQP29nBH5nGcko01dmFy2PivXO8+88pr08/n+PFV8xJ+lP1
9s4+YhfI4nV+YMZwJAVkvmR7mhFDryD+kH7zlZYG8Rcf4AljOKH+BfmuhGstihNq6NUWz1TkUX9F
3AlEKFZ6ne9aiA7BcRY9JpWW9n9uJD+auFSRYlm6itA3bFgvFmcRD+XOI+J27Vk62Is6Zw9DqODu
fx4FSt40o08MNNI6/kdABk5gcx/grb7azl41RL5xokNk9RTH//e3XwjoRS60Ell8SHCVzfxU2nGF
ifyBtnMVHEVqgpAVvubrhGBK5Q//ln6Np2S6FdHn9vl5PV1ulXu/uHpgFbrj2GfD4hCbnH//K+wI
jpaWY7czWQikP205ssSQXKpwNGZgz+7w07yFpxZQhOBh53PpetVe9fPX2ijRtnTGidFq3So977nM
abgJxS1JgBPFC2M/LIMnBe6GW4lEz5zrrg5+flwnICKXaGfwXh4EtYKR0v9u3d1EKECkbXj9ip2H
fYhSz9WIBeLUe1C9fr4Q+gGSxzw0AxYhoCv8CWvKtkxzT3SLoxILM/2VW2fvl3TapgY+/CKsMwMb
7PTytv12Jbgmsy+K+QBZa5Mx8GDuImzVMaoIQXCHhIjtafKQ0SOGHWeGhiMQQhEBbKvM7uF9lU14
1y2M6KHHXuGCHpsW2egoDX8Z2PYpQ2CSOmhaUbT198KhL2ux87kYKxNIib61uw+iZf449il7cogy
NQWkuNbDZvqp7sxR7+CYTGwt56z2sOByRDsvy4qMZytW+RciXnWDMb/3hzrk8IaZMMYnbaqbkvgG
gUytsmrEd7eqWGrBVpT1PMCb/Neeb9pKkV1YpkGG2FAODp/cxiBmqncUs6KwuX9RJfYfzoMZTX0T
kWZnq6FcknpNeK7p6ApjAdyarCtzl1UsoHFlAq1sVgSKxOoUuxTe92EYXZcqYSRvkqCb9B+GoTR9
gfS5iZGBGGLwM3yCScxVV5BjzhN0XnV1SN+ECyrMREgAi3FntzUqeGUTexzhLCQe34ZffSoN+RZm
PXsA1OoG9EBr6rZrFsmlei32Zme/qSjTzcHd6UG6f7OxpcyoE1g4nBAd/1uFce97WprOMWls57O+
v405nQwZpYRHmJp5C9DjRA87KBx9fubKH4h/2X9U4kmMEBrvfBWcJTigLG/t8uWymENCRl2p86pW
t0qEqtmQPsiMBGdI6akHaKpsJWzYPQP4gmmbKj7Dxsmd49M8MHkskXD/Sak4YEXCojYvKH7lYMkk
/d8lbzwJfTR7sEyoYFA92jBa+aABEwjvJerU72IySaKCpcJaaJwAE77fiby3TOzpWBr//5BBDMww
LJEHoxy2dn8hcNv3ClfDOeACzyDRiuI/ysIzpFk++auvXTbFgSUDRNzSK7a2FgrnRM6tlhLA6YzF
BwmoeEat4AVQ93Tbxr1WcS0jmuOgytTSOmPwo4vktqp6Nfcm2QeJQzgSgRBjRwLCMMawRs141Pvt
ZNsSpaFcUDhS6BHcu/4oPSDuNwNYd1gzCIV5sRBnwphfpSgIntLKa3grGOcicaL8AUlG8NHtsnSn
2A2Z5OwtwerlS+IRG+2aAZH7EQkLeHz9Nk7GCJAibIKk3sQrt/c2ASjlfUNFTgiXVlGWQZJHeTJ2
dy0j74U+yvEW/DHscGBMPKqmsKChS+oQ6tQayfpimJDrPUqrMTgn0JnV5S6EWW8PPI8Ro2lQOGL2
LyhmBWGCVpOkdCrTVr6tMvZo3IrOwDyCSeLxBe1RAh6edITX4DEg+16LAOT2jKlGk90/vQXM2LMW
RAg7Z7vvPSHj0zUsRSU096HsZtJYsVCObuzqICK8h8wlPhpEaDkZC62q0j1s8S52SqQQJEP2jRVJ
rSqruQRTEEewx9cCSTk2XpVzmyHLSMerxG0pSJNZNikiLVziICf4o58qzJnIoayuUS/p8HJe9puf
ABvylCL0N/n2i2RHpaYpIB1N+xmlyVs7aTFP9PlLCDEEr4KKYggDtJNCJIm2YdHoCtZRVOtVIDjC
x6zK5v5AR0tPtiv1k5/bqL3utSexY/81IBgD438RAaIcULKIB9+zZT2/5b4Iq69R0WaiwHYnbH/p
kpCwZ21y9cjQKT/TtAxW2hWg6eqBanaZJUj/2NECzgB1cD3RQGU5w60kP51MDEg7OcpiUrQZ+62L
O87SBIDdOk/I58A7Gc1HGEvC8gy+mDiQ6La19eORKF2Em8xFHJR7M0tAJ2H6Fgpal5uMcYUeWnxQ
wgZ7ru7OezmaCM+zyCy5Ib9YdrKbPH0kqsG9kFY/jkZloVlhVPKGslzDjVHGLoT0tVlc8sT7EIOI
T5m5XHh1tfBZaXVW5FvOMX3rDlLB091fAY02bF8d4ee2CsHIH+lNdOeArROIggwoIYp+Ik4z/p/c
6a0dbVQVbbpPwE25GPwvjcgzfru5zSwCW1lpHMUmfcx8ttZ79aZRR8TjEkefHT0BJqHjXtohwIoq
5SCM1PJU4K16Lz1+rbQDp8gr9D0sMOI7B1xTciK8QN3p9/zH8VTfiQA3ta+zfydeWqUE46upImb/
EeNDb5k8sqYU744bzys8rgih3bIqJzQh35L5sm/DQioNR0ccbe9cW1Z8T3dN3ZSruFmApvDuYIsi
dOOmi1pTtOt/ET0vlET9PKUgxHEVbn60VpSmPUyMaoxoXyuW9NTIfiguFTES/k4UtLrr4Qe7N6Ek
pZM9aPSITsAk0FLrNf8oeYuX0ODCoXvi/i9Zku/UQmHtzN5cKRqG40TzRbohwh4c5tcKODuNmw9h
rd33ZKrsHeLGD1+JOwSaW86GAevd20GpM0rC3tk5mZQ6w/CI+5NmGm59w8iEwICQFwkdwfX34fGo
DgW+O+5KJm4+GOS/oXXBIiUkXuJvYkg8K5KHkP+1uboilPkq9SdvOOTG3r37a0ybNL5SeQHxLNkd
8rpWOr9OVHvsp+5MBNupXW3wtiAskUdZGnlz2bEvApConOSEb3OWs7/VWvcOl+V5UWHvCFsq4X39
acSyan9LjEcdOatmCH2m6GlWROqmBHr5Dtnt7z0xp3KNWJXuw1BBwQWtOgNvMCB2y2iDiFJ3RKTH
LXOJdjtnUrpWPtHl1F0GJPsv46zM4ljEtKTwsnJ003oO1dmnMxPudxLMPk0NClXycXpFpT6+mYUU
WVwpeQ7MeAu4rklGbfrgBlE4tpDgFXV2Bd1phRyBKBRT9aWXkeiVM8bfrCF5yw+/T28nJBv13YQ3
LGgb7fxUGceMf42feXk1L0eF6UqQw1FX92G3hneYmCmLzLSkTPOLJge21UdRCv3htzrpyg9xjzr2
il0FOgSGAcdliD9oXN3q6dUS/9YRrrT+afLyFZt2T6rBYU2LfqtFhliLpIeaAyqGI8KsrD7YZYkD
vudEAPBvpgZdElaa7R57kZ6hQd1aSlzm0hF0FAA8NBB46uvDNu8zZDb1ZbokKPRxq7Jbaz7+7mWV
8WlKsNucInkeYKC7tdxAGnKnHLhqRw/hKZpqhiftzF+Qa1SA0tKzgoMzh9ZQjM9a5ifwYDFlfKd0
JhgGEs1/msGnvoeD5J1ktt/ATY0giyvVDUyuOoqpVhImnInaPvX8DDGj5XyiXzBI4rap+uhTyEZL
mIbgmP6K6K0gMkWOH1InfSoZnK9xrkJniMmTV/7QD6ha0+Y7zNayM++21GuJhVq9EAq6CLn6+zn2
OARSaO0JEdmJxEFi4R8T5wfxDfz45T1Ue0cHGnhp0m0hsLAwXP8BnVMkTjnCp97gHDmByXjDcHkQ
Dt6+ZbI/XYql9UzekB5PYuuJOIybC5Cl622ThJlJcs7+HNJgKs9FTOMVntDl94/UNSKc7dLvDbJ9
tM7xkbdZRtbCo4Fn6nAMPXsCKEJ7jxoi3SaDSBu6tw2rIZVo7PcDviSZfHuAaZmlWPL3V8ZP1pu2
g3KGS+TFTJWZU8jlrp4zOyjA+VNCtI5uJXw3pFigg2c9Yg1TDsrXlBHG/X2zafXILNWAEb1FQ3lb
CiHh/S0VSMGUqmKKFi2DnF5NvF6WGqYX++mWez9rpQq5kaS9yMmQ8N1MPeGazzMQ7Szb3mgvycDg
U9ha7XvierL6pa5IwsVfDfBvd7iGZhR0Z+xQaTORlYdQ4s3PiVoHP08Zci/NufaYumVgFASTgO8i
yIS7KRniNWfFYjja1EjZRgTVWQgd/4zRBR4yTKQ6z74BWo/di7/vRCreL2A/eJlqIin9QTfCvrsc
75CxPN5NcjOHt8z928yh7z6UmFOIyBVUcnOIuaMwvrQcx5JWurcaPOyvEEHz5KHjRJ2btPmf/Vlp
9yzIWtuOQf1r4Iuk+0QaR6aNGYFj3By8pW8xThhHhXHUWwbgI9AdH83aLpcw37/P9mpVOEjhToZ/
ByoJm4IgfTovoLHdh8xb2HEXSeJaO15ro1dtBO7WnzsU3juqOmANOYXkDobcyCNkRYeMrGndzA6V
XEKIC/cJIDD/1QqeWMco4dWsyLkYZBKZpmPmHSaAIdfngP2IiE28oJ+xFNjPPQ1bnlQWFXwiujo6
gWtosyXzWV7eSov1AueyWdoj1/PKTDKStSdGjDfZSK5qphj+rL4cqb89AX/ZDcZQQ3GzDXCXiN1/
uJkt1LZLh5TFpp3O0WZ0Ne/4cV0NoekLSAmaUsFa5I6rv59pDHxYAN7jgig8g6YlwBXQPd3Orh9q
sSWGzGGdRa0Q8xZfm0N+CMBXzL6YgzkqmGRGhr6EO5L1pwk0YE2qimXu9OmrWxpResBReqQQkNSB
aLKGBk1KE+1czgJ73bRjbXw2dK4/IjV2usWvOE218YjSzp5nX4DglISR/CXWn6CnnQ4rD12L74Nt
mRxmj40UAOBw89ImAS31T8H5C0A2HuPxzaac/05uPkSHTrFQcQ2Q7iLvOJxcqx9sEpZ9og9oL8Of
qIzxHF0RhvTXHY0XVL7v8brUkwbbkSBOk3zyWg7rbpar/5iGNOGxTqJosuqTCy6SNJU5LvgZRK4V
26c83fh3v+YlyZzoec1h8hscZbuMrNFKM1+7Gubc9u6z2Q1+89m3M6B1hkXQYm6mfh8R3NiO4QUI
sCzDnoMBmjdM82vWt/WPmpNx47d5jpY65G1fm5P53ovjxWLXFl8JRRgYPv6C4nFD0LTuqkBTVaQs
XzJ3fUeb2o8Zc5aLY7YQhyZqgMmL9fC96rd1P63KeIfw8Yj8NMMQSkSqrkq1Ye/5q88DnJc+uemJ
E8O2+wDbWwj34lQs+NUpld9FBBSaRhk3Hk1y2y7XLoU/OvlJ0zgqkGwdOTQBWlmxLP6x7yn0NsSw
pJi6LFe08lUloNFZqua73ZsSS1nu+ljmBgsCJtwOXPsigdA+cXZ8t6RXvjdUhWubG4mYsECieNQW
rrJvG2KNvlOFxFpQAqjgEs7FIklLohSCFVHKcWanXlTBDh4TIK8EfupCBQE5DIQC31k9dt5lcu2J
aDE5yeddDD07kkV6RRC70s/Lahw+bOSFV6/vA1Wa8VpaOLUAT705MilDy1Ci5YyHi8Nem8Mm9ZQx
Q1v/t9VnXVP4HL8qADoUqWNYKSsOMgCvexG8TSCVtP6oZHX8YB3u75B/Hukewis7TgZVhINmJlXv
nRqFUTgZpR3/gbZeQkPXFjz7+XSz06KByumC4qEaanHoZfLU2Mt+tuGp0acc8dQFyOAgX6TH7A6a
iaEtvbS0rDbbmhBf67OZUFbDp1b4fM9E9TuWcBfwyp7xU0ylzI1pP7e5jK9gcCFARczgdg8rbMS6
y9bHSnLvQm480B/nVOoA2jUd7V+UJbw5QENnvyTtZC1R3MRisoGrUiRxU6AMOULhGnDlHTFZIG8b
VdCBx3gqXAjqUwRHxthCFo00tBVA2nCOWjCGIi8pZ2OiWRmOlj8D24uTG+LNmQpBMH7nch67EWOq
g5phEVLsfubhPjxvJklAeVPi0J3jcx3sMrVMP9Mrqm9VNrQtV3VtoZeJtyFHjsA0vmDWtRuXEpzG
JptqA3xdpoc8sDaV2/LBkm8KH7Qf7zQjLyhBnbrbM2ZRMDdlI5hsFUrZyjplKs1ZzjNRHWMrfkos
40IQq80zAtax8PP2AUKUThnVhLWpdTsk8a/R49YcznlYvKDc8Z1k3uNThH2o42jTk5xVg+cOgJO7
Las65L7ifN0IeEBYrc7pI8k97+Bpi9rDaoVp8SLVh3LGreXgg4VCzePt32kXGDnykYTxm5uLo1wL
uWiAKaP+M5FzbJ/Ah7LOT0R0yr5izpTU0xnb+0V4KgRdz9q+tngEthn6gLQtLlEENT+Z/IjBsuzs
v94jmnupJO1uA6WzwVKg4/3l7cHWO7qc6OEw0lMNwvJARp+cVSf/8qwSKJmL4lFAXmIp9A5QbY3e
Jzm2ohLDCOumM3cBfV00etb13xQ9KesrHlqgbRAcg9QVbCfQD80c24mGk9YwLGdYJnXst+TA8+1i
C6UDQghaUw92xLH6D0oenPgnvKemHIiE+oNK14RfuyEzrxwhi7WvPmYmSboVRlNkETt/l0lttOul
iyCWSY7c/mcQCHjs+Hp55ofx6E0i4feCwIhX1/oA10myFic3BHNjnxGpWbI6KTwUhfSxB/m4eyPA
jb1/T9BED6tp9wWaNnSiHtfJIrGTlsK9EiaAOdfA4xu8gxlHq1jh4yX01hOKxdoemNM6X+OxQ5H/
h8QwOOCGSnOt3rqARL+UXwFMmL25+Lt616oBGObHl54wsTUGDT0Kh+hU0w0WI0UJHADfqOg9OCOe
6XoUnvBLRQ19NgA7eMA+EBxuqo4ioA5KdCrd27UReq6MpWeHNA/VCZ70mJ2JuoKD+oszf1iegUVQ
93QtyyJbxMcPwpCJGFZY7oQX160Ctb64fDE2gI9r3Ep1tcLHpu6flTX5C8PxWuDP9VYrUYX4oNNj
NQh5F9bK5El06dN4D9HNt2h98APT8ELb0mQdX5sdKW8m7alq3AKzfDj3eF8hTEoVZR0lW6JQjiS+
5knS8NqN6I37eDTLgi/qqPYhE/ftlozzmABnuLd1oGryrrThiNAjuYgX/QkCvL091wZw8tuY4XQr
B7F3aI0Sx8nYxQ6gNz2Xnj7SGVxbRl7kGmQ8nDtFbaeTDq0pemLYqtb8Fzibb2b2Ts1JUy/Ajtsf
mwSiGd1jidRuDpBMCpN5zGODotS5uKCdCfT30qd74o1jXMUwxBiMKtKbOjxJhcQS2hkmQ/uytz5D
JCapj2QV8v0enNH0FVqdvTu5eCOqWZ60XiYI5sH2EC0vd5BK3c6UpIW7Oa1NxfhaB/hS2arIS8eA
SW+d5aGmSkLPGjwfsLPw5zrfvx8X+oXSUaXE1/BEc7S/cIaBmSN7KRAXvsRs9gQXVEw5rTJ6KiM7
iN0lIg7PEwa++ThcM7pZ33YCZ1GhXrBqWW7IJS7zQOCoQ7U5q5kTGO74JwFtbpqG+Ihvq0Oo5rWV
GBoLJoi29XckdyHTTTR5sBt3SZ9b8DRr9jgjcYvavyh2Mwss0oZ2ylZ61bjuhkQjfRqzKNtTWQAl
e22xU3DVj1g9MXxH5Umpa5P+OtVPmrCEvIruL2soygqAR+/RdZh35a1xxaudw6YVeBjYYOA++nht
4t8XSnBf3AaVllPY5xuGm8v0WTdJO509epYuR9B1/YEbWZ1L1tSDQWNxRUe8tSDYFJti0MAeZXwW
GPmZndwREAUbVYMKB3v3vP0clmqYdGB818WiaumC+5VVJ24VHcLgbddyp+9SZJ5FbW44UuD9Uoyj
aCN+TJVYNGfSB+LrYWzNc50AgLA4YUMthDBZSVTErbS2PSGjLYTdGy5bRed6dgjqe3Yrjddq88I3
p1ZUPGejGsTZ6H9t+gO1qmyeWgvuX8rimxwi155PLhg+zlhEi3y8dzCbnOB1pPllstJvch2QiT0a
X7591gBCHN8y30ul93oXe/1fkZUsZcnnxoS66++TXzt8mByZlaYQgL7vHUQSF6GLucm7ox2YKr8K
/8hIwedvDFOCen2Jyziydx2PIruyRbEG7g8g0xRETZ1t084iN98TlE3TcprcO34mEMNNi9gLTUJA
nWIxv5EdtHKaa0vVJrz/qh3SkTe64m0o8p+Yu6ofmaQzt6ame9PcUoQzkZzuxAg7V4lh0CQF6+bd
GMM2CNP3CfaxF0MFrKeYSkSkdW8qB9d6WR9PrYrPh7lYcx9O8a0C/yOxxH/y0j3mH3DkSVsw22iN
G+isQOjwu5lmUR2eTcnPs/Rcf1F226gue401jR1yNOOO8SXud+Mfph6MXkVBgzfr1sK/Sgr3I4/0
xVmDCgUeGIzWTVDSpME5Lpf0gUrHExxacXXsG7Fw
`protect end_protected
