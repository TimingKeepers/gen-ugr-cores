`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SCUop9gzf4hg+dmpEMyi+zbT1gxVfbGAu4ZGhQFZy5njnFOjmnZFi+sUcLh+Oo+Q7FX4ihQduxqn
tyhEwQ4tw7kdoDcgw/PVTQLaYj78yjl8aBG6TDYW6y+2VhUyixIrdL6Twr8RLDmDCkJ3dEdBMteD
DeF3eDExrpL1mIKIep8fQVU7nACG5Idqs7pX8jjViLCQ2Fz1leYh+R9qhuyIkpMyVZfOM1FTUvR/
JVHFa+PG9phoSsO61D6/o+F2JyvW4/fSQE/ArIBFxKqkGeFEKMSfhW0XhZiz8Bo0XILVKk/Xhx9l
JtcM3cURynHfk7LtugM9fStpCfZcg4ym5+dwqQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mz7G/IwpqKZUtRa7t/axGLKpNWLNProYsC5mKTZgt4Qxsm892JdoUXaE9Bbe9BQ5640kKsP/LBy/
lV+HR5RBo4i7Air5k7lxrCDBSZgZ4KxNhal7eNEGYex7c517cQZrRRLztS/KXcX7+NDcm7ZwtOWV
fDbfnYG7IMmbcGvD51k=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
S+em6x0QxfE5KpieoXm2e1zcq9XpaaOaHVp3wEg2VlZjHupOwuwxjKJSgYvySTlCCCW70J7XPjGz
VZ/VQ4BAJaeF6yh2xfGJDNG6qahqqUvrgj97juCE08Yh06vCYUMNA33U/d9awPkii24rVrgLGkYc
FRB83/HjhQpX+a5LNCQ=

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6432)
`protect data_block
S15aZajJ/SnWdqU5nCYXAiH/m97c5MLVe6k2l7XzLbg3fr7vC6NSz9oEMTdJjVwLBZfbzzW+NyAT
+DCGM+dBw1Aok73JeeoI26NFnqbWKaEPLG3qdv5BHBvgp1z8V4jFMkIi27mwrPbpm5E5HELe+hkV
CHeNyABJTWtwyOtUE80wYek/T6kVs61dYq6/azK5fNkwSJSyngKSBp9tEkfaZc32MH84Bf+Ojkya
TXJ4gSpiPfpsmHYfQeUDrtjlRXUmPEZERqOHnVG1/PhtG6W35TAXGMcLEfJMegd7NTTheloa6E+Q
ZlNXelxPF+SUxQdJDzc0vheCmCRKRDaY+vsMKk53afte/AEML23mQ6jR7FzklRsM16XfGEPoa6N7
tLZYLaLCaWgA+FaiH7+s3ZxRlgAGOQGcjwMOGc2PvfuQcTaudPoz+OVGqFKz/EZTLjEzfSf9hVzM
zPmUfU+zir0jQ+4SUiSYAmlRSzNvX0Q7rvbaW2knZEiEgqOfkJBatZDeoTWwU5gGtR1qm4AZGS4F
vPxqlhnC/IJmvoGxzGqsjxb8sDns1xS7bdN7gG9rd1DnKwcemKiInW1qe68zs9jYQ6Bfclhrm77Z
0EbLB2NhG+QY7IOHVhOnJZ/Pg5BJ5MHmfuyZ8HWCSZJoak2u6q1RsUuAGGaduSLmn3FFGqqjWE2Y
rU8OFri0AzYkgi6+OnHP+82qkjM+xlHlJFRRYo53Qu/dQTbuiManHTspVBg5BCNmkhWgFpZtei7k
9U3t2js0AhtJIx53Kzf35v842b8Ll5sdDmuh0x6i0KeTffLrL9QI5uCNsbp0PRTIkqvOcgaLcGgv
U5414ud4BfPGcTphHMycMi/2bMmxWG3QU5CfwytntkNpLiRUXxltuHIr82WrlhNQvk14kSA54k3T
HGn80Qv1Qz/FTbG2v0ttAqFbP8eI4CbguyLotFjTjWJCe/LKUiMccRYQjjVE3HR9Z7vFipmuWs/Z
ago+arBBkd+XukcsKPMh5dq8frGGFVIW3U3EqNOKRyh4nBhCMBa1SlvEHjfk8nzYm5wg098wn1tM
3ASoZH0N6clC7lLNKBQgO9FDlKlaptwqT1mv04gTxMpnJ3z4j8qJFxxtLS3WZTRszPrJxBNo78mb
pAiI0LJWb88AAHUCTVNqN7bhTM9KIOq3abzfc8mPYil2G8AFsF720O8mJovImvfcvTsP76S8JTDh
m8lN1rqgnie4k04yuWpk8SZa4CP4dLrlxXxhRKUNd+ATTIotSruRHga/X0mXHn8Z4zmoWK/1QL2S
3/1MIVImatPkJGYwjQNwmnxTIIayijoS5RTUAmRb2VoAoGoBNaBxMF4HT9XAMOErSMb9rVq6vjHH
+Cbd1uEBpJBIZbpSIusBj0xYIrs89Hfk/LengpHzPGFSvKq/1DZBQ4Acym5FgF8XBPTDkDAJDssK
bhPSfn2R0aFujiZrWKeLk6wqQ98zyp07wD2eMSstb3jNSXLUmR306JXv/R6ppjGe2FfZoYnzmjRS
4CG6q3JgVdrET8qRqObInVs+Z7RwGZUYelUYt/ReozO5T1jXpvRk5O+h0e3iaOV4U16Z2FFISC+3
FPHv7t0fgLnjBFQOC1xxzdj0AQU9GrUKHCgndHUktu6CdDwjFyfgxg/PFFlHU2qYw8UGYLnGURF5
lZNixFNRo1e9cfPIDDfpRurCL1CV31+5yz2A0adhDUa5BMRxndSqpwhAMd/16x0rg/PEhBGZH3my
Xv8dsqYO48NDNmsQgpOh9FkaSs7x/+oM9IyF0vyahfNA8JDjhIEqbIGTbL8xUOtza1oc3GhmW8Zl
QrpvQNR8zQIbzvzamWaeH4TIVln5ZihH9SsvYMqseLYtJ1ZhkjmnPbVHf3/IoNsE0DVWJHNX/9vT
YCo3rh+4SvdvJi0X2cM4RgyvzCbQy+RtT/5eaTCnxQC7yCWo7AKg/SyG/WDtOcohh+51/lbKy7yk
k6kFBGdjjwF19wHENtvtbClUkkCSRtciP/Ec5/nPGVTgrjGAdNAo3pSSgwYbFzbJH9fbded78KeJ
c8DTX2HFsGB2yTNLjFmTwh1/YQERL1RSMNxkLKiT27bSuRgBOVAXW8rdqi6jb57F096KEA3v9F1T
QFl14DA7d2iVUJRAv84CxdZciYX2fToYVAUiW3obLMHI9MOBE7ET4bpiwucD4ZF1W/UbaoUKZpdk
CKM0Ayglpca6eWsux/LvnkOOBoGefxJU1tpy1rkzzhVcWLXGmM1KVI8J8BqNPJUobsvPniMYVghn
tLqxPUNQRzrWt35WKGmB70ZaVuyvLi9fuAJ2IcFPD7ie+7FnGbaNQHAFeGnbdhCfzjf2NwLz/oOB
OadH9HM1D2koJh7tlpuXOuMdyI9H1X2CFV3A4Q+8COWiv6maoCo/KKOuV/SfCYMmOtE0fn7D2Qcn
3mKFokO2RwiNRX5ph3UkOY/Im9rtCQvhNaEDAJp+/8l2OgGNB5BCWg5PeSD6OEDF944CZVGuHNp5
VNflJtBNvClxubLwS+rgZIeJPo/gLZ7b2z/didmU+kw1M+US1nPmNHZCLeBtDem3WF4U0wzm4f8I
bVdfMgMhk5jkJ7DaYZ52wjuI9l1pIEwQdaMK84AI9BGoI3yY86JWHz4ttXA/OQHO+S8dRqYXGmd+
MOWqxCXKcJM2VGywLFuEZtDFJRkN95ZhSKqa81ZyaCDqHMrZwPPZWUxSPl5R48p2xztGxKC+Vp8n
rEMV2NQ9NKLxgzWcCysAxdkm+EsL+Ydd3wfc8hRTFq5i9ptRYC4PnaOe+rin39VXjkQFDoKblBIj
QFQ8dA1Ob9veY3ZwyKCyK4IsQpCdZ8/V+0/Z4RIlXosRUbiGoi7b5MQZLIhzZS/SFwI2G2oKJGzw
sUHpDE7w69kAU2+1MSWyUNX3rj36z3iUnYQG3h1CZPzuYCzG8cSxpcEr4XQZZmyOtGgxa0G8qzEr
865Ma4uyi/glxxVs4rQntzBdEbif1+EaFfwA/j/eidNDtvzepEgVlcl9J+YvwY7I4O8Bj9dPYhGP
asIBlnoSvpaJNAVQgwaXSV31oCMh/V3XIR89YTIM9qxcwL1SEdiS8dpzlrr1zq34Y3hg8+A0bDZ9
4A+fElFDcN/fydBcXtjqv0WVVc9S+2rDgj4QlPMyY1Ga8x2lw/Qqks/OPEOvyZIuRzab95KXBPIc
ILXJcUHYqmqqeW/wOBgyypsXGtkl4znedTeyR76U6nZ4GC1eAk2i5qZH8+mTf7Zb42/ox9VUIT1p
Zw+vSRIz3hrQ7EfFf0W/Cgn9OqYpN9ZXoykSERNtbD6uBfrztimjmFNJKcdo9umTEWWNgRC1mBdU
NhObsldAS0MAU5D/SBdnOAEFvT4CNJwjiDGzQYEB0UkdgPaE5CBu7F2dv/HXWcf5ozLnDIl9MRA0
mtEqZc7hGbd4EPMiFI4IAcQcImT0YYtDKuJKQMOUgdD1DDqAvmHK+WsZIvE+0OY4U74Ylx/mR7yf
PJXYbJceG1tcQMIgvwbZb3d2yIxWvq5rUrjB4pBGpVEE3Ng6D6Hw+YUJ415/chCC8CDTav1QtbvF
F9hgmSvlCeJ2t1JQs0TSEnVFuUzk3uR3OMJKH92NMfuwDUODuN1R/RD8GwEwJgoNRd6NCx63S2Wo
giNypSZDC7SIecknOO+ulgimzkPxXcHw88MnPLK/XgxEPoxVS66JqyAwkSPdhUP9SjRwB7UkTgQV
7pQWSKOw+MxjU2Xizblh41dU/EaBRmFKmDjv3jF3Lhmy6At80r1e/5rOdkZswmfFPlW+nS6pJ+DA
inGmm+8dCRdcRXFZx2GoMtE/EuGvS/AcqqJ4cM6WqljoXNtZtzaOzBvjI6aCV1z2gYKRftYngtH1
3vWbBkvZvIsFoUQCL2CyTYm3fAkqcn/kNhyOsl+nHuzHkzVXp7gvwcsOBmAURqCmQi5WBRzW3raU
1yBxMSH7iXGFuAcH0re4RuVGkFh3XWG6kgVUeB+BD/sPF8dusYQ69LG67e8Hys7Q8izejjAIXoM8
rBQRSf2nJZBy5JUeTmz+YMQjhymIICHFEdJR6w9jq5fPRwAkvaqSY2N0jAMPf4P5wn709QghuqmX
T+6mO1XrEebLg5f9YBsd0uwrSSqLlr6ru+EZhZXbTR8PhWbuYRLna4ZUzmXl55gqGMse92U1DnB0
dYeJ986b3LLcDXjxUmEQamQIR7KA9SvL7WAoGffj0Y2vMKFhxx8B4CWMgdIvxqRCiA+eKoepDpPg
QsaTX9FYEXpgc8p1RW6XNK/EnNr6zAexC6YuNzj57frzpWhfQvKRYD4I1aEwTxBzGFIP5h1l4sLT
jtsFi4OuR5kO9676AvAY0JiO8z2HC6PC4ZJNGU+3kKMHw+kTlFxMJKmvj2Q0yrgmTNYxIjL1w+M6
2KcSVj8hL42kI4Mf46n+su8iSBQgwkpE79ujtUtY97be6gHH6C5MTEyJIl0cTxfTKDNpO8+iz76x
ZhK+kSuiAS4+uHpBOPlfEf+5uwo72DVnaK3zno3NlxEbzs5T4qmhCiamHNZfnVUNwFRqxv/roLy+
S43/D7QVJTzvf4ZOXp/PUxTPIK0v/tYK93UBBTr/DFkiqADmu4vC8HrVzAdo+VH9P4y60S8gAywF
4kdF3/morZW4XxiUCBVN9sugTTBAfFfoU+2C9Dl+5SmUpBtYf9ceTl2QHXp/w5XdzF3qde0VQBgW
rJhVZdMS0kcpGDKd/rp85xB9FTdeOqHHqo1VErTERxVuDrfYrwZv37lK9/gtmkok3naUrsJEBD+s
XCWGENWGc0S6ifdigKDinTmaNlE3RDd0J3zgWP1qhWeipR6+RZs/thNcFj1PvZSfXCP+3ZaMbtpO
mlpTqcKy2yiJCDAI19p1YfbTY/GbN/fCJTF8XIgkbqIws24e+YGnciS/UyKFPg1nRdxYz0X+5s03
TWJyd1WYFV5sKSCUFz2uquubxbG5UeoVCmp6JbKtO6bgRrALg5+WpBieQJvPk865FAFxLgVvGCWZ
gRXWuHfskMdWWJ0cClsq4QqPbSyrO5Fdjo0+n7re4MbgRd39upRVuEYe7IVI8L+Hkh1+nEtWbpLo
A4rG9wy7Q5pU/kWf0P0x2/QrAvhTgSxSNfvaVLP22Wbrl/qbdmeJ+h86nvPZoI3rPHvAnwFBTzzJ
ckT2XdxUwyJ+zxRrKBu2CuquLWgOD6SIt4LyL7MgBW5XBBZOUAODtKful7HtUsCTdIfDlB1OZMWq
CPNr4JSvHn5Kw+3cnRJkASYoViIjPzqjptSMCGr59l2RMC1Z/ixspgGod/a2xMYB/UVYW+Hipx/v
t22LnzQZxZ8lqF0Y9wKv1CvMHsunq0EthQ05fzrHyxG4a2D0VHiL6xz4sQNqPKDnnbD4me/DbrVV
UVBr0PqTwac3FAqPsvoByHAyfJ3iN3mBWQ5iRSKqG9L4SQQ8W+9Az/Dl2btCYbJR/c8mqBwg1Tzk
oPavBQadaKIkm90pnyk20WkFIADBrQnBlH2QVvKlcYKtGgBqGiGwLcaG9OeDm3dCZspUDRfycYQn
Eyn3WfQLGnhzzkFzJsfrTI0oEEyB/kak1yfys9Gu0oBKyYSKQecyz9xW6lgXYzKVdyCwoOd4vYcF
kA0HEfRoQu7geZS8Evpc1B5MxLlmOUTEF0Q6rl73qZWA/ooMqht694Ak5UBLZX5/amaYK5yHWgjp
YPzFVrXUxeR5W/LiCaTbIcoyV23B6Y6V68XF15cEzMNdgf8XChlSerTuS5rkO4g0Bx9ApKZdMhJK
u6PMWu0g7JDerwNMWAFs3kmyGHpifGcqQDNDuo0VfgCGBx9Vv++Hk5GvhP0eA0BG8tjHFI4+wpfK
zP+UXHG9KvmF601a9wJ01KsLe5jXBe1r9DHnEbqQYL0/fCeju/MmG57QSBagLwXkHupIzMIRSPyE
clD7UiGPaOd8zf4EQw18eRmbb2qGmlg6odP5q7QUxZV7GyFb1iqiqprfo/YqONKP4gUR9bMJxMwR
fbqNRQ+HbqKwe+tdN3Bo2/XMFxRT08rYFeqBl7kfrVRyJt2PlaL18/jo4enD4E8RG0A+PIc835gL
k98xKlE8t9ya9vZGyedkrvYCezRvRajIGdc+spbcEaAXp5FKNQJn8+X7omNzguDy6CaPGbI4HJxB
plGuXAgUfr/Oae7o0l8WHtNA9vlF3j+/7gpyj/WQSOTLo391J6l5cMsM+bdADnJuLDV7lohzQQDs
+8YnEEBz/QFYguksDhQ0GBu8d2QUpgHITXLfFtR0TeyMeeQSPPX9JhW1su856IUQhsV872E9L6tA
kF2xucEH4dCv2nsz/ut8E9ZMfkYKOoUK2LZbbdfrrSLih4p7O0iMmblyCPWLK7B2Isw5yYIb8JKR
TSB9NfWMf4yR+Xi86/R1AI/4OkiLf7wKkOWsYjSrdQFy7728bolaMLH//IYbS9NbkTU2Df7T8O8S
SWf+kT/alLZTuBYQgqvaVUpU/bUIaCL2XL4Agl8TUNziCT1i3leTv+RMzR4JI/MfH80mmCSE4KmW
l8qsD7md9EmojgiNy0jEvYbpoEuElou/Rpni8mkaF8DVGnPgrkKQ8p1UAioPntuYDAMloPC1XUSV
kQlvf59sZD8V38opz8WSR2zIEfHrXJJlWLvdvLVTcq3qIVkfF6w2FBcuSzhprWHTspPhr1ynh1gI
iHMXhiGhb+s1zdGmHq4uKSQe8GUW7uQ6hgJoqSgEfD7hNT7odMKoxmZwILCoSQQbTN1YBd9AoI5n
foZ9ju9eqN77dkCHtkX/pMRyE/SsXZGnQonXz9wp2hVKvXot6SWgs49Qoi5EzPcgeJPNW1Tciftf
qv25hzL46dYoe4bvTnAO7H60O6VYjj9U1WcD/Lspm0IndXgq++N6jA2eRdd1usZlmKtGw5/Fr6r8
zyzecMT2Z5RnIbudF27EXnkfhozk99UYYTqmAGObsByjhMpThEpfIRc79gEQNQj8IODEOsUDhXJY
ew/x10GPr8I58grxeVycu3/KkVfLh2U+7HoVWYIaCIg+62aHY2gVIuGj1PHoixJEyXZn6YSxsXvc
MucnTYJxaNNXRzx5jJEzu3dtF2+GYbLpWzBB14aZ2kKD7wRAqQvWcKsFsBiNboW6Z9+ISnXEcA1p
WUaPvJhdXGugyaKjzdgN35+4Z47QQ/O3iUStEF3Wd3QFfJ0iYGU1SAiZUcGBffx50QfMCRclZrQR
INO6fuHdVhs8us/VY5/ITHD9bVa/jyvTE174ottf1r6RoxyYyVZ3cS95MBjZasxyDWX1lyVOr8TF
HJO7QbNGZBPHj2CghJsaDjqhifG4BsbjAbRRtQsoCMd8zroDyptSTJpM9GEC8NC4v1MVxTfE+Xkd
TiV08paWzuY7KKtZqi0ivqGmfrkF65WW4n7j9betMtywkVMUD4qChsCiMRVURgh3/a4+UKAdzFyl
7hCY7d086Z8Dd/VuTBz+PreH1ifNChXg0S6omd6ThMiZwscgyED9lSKQXfz0B0HP1NVJf8r08H5i
6XJXSQ4eD9bGuaxmvzmFEDmqcCyaco5mHQDPGylYA9nCB6PwI03N5Gkp7QJhvL9DrdyTn/UCWM1C
kKtBlrbX5aqDAmFVVzw1VPyBBsfL8dNgiVK56EjMpk683ecQlxPKc2tZ5AtZePFPflylB+R3mR56
CW84SuGftP7MnZMGDvFGU9izpP5DDm247I6RybEKUTirRvkT1CT0ucbI5t++B+W4V1JClAnKtv4i
ayuyLWl56vdoGpDjR9O1tqxqj7bKQDU0qqcdIXvG7+bACNbRnKmH5YeAYWqdvis/8q2Bfapj3f4J
+XAW+gxnp5pKnVdsL+s/gGMH/dyT0dRYc39QvejBNbmJKXl+PGvxNwbgRbP0hvma+ZPHWVhumXNx
Q2c12QeQx08SLmPtuvPJY69B9YsOKhHOHL0nC7brN5DO/ioqwe8hY/Lf33HUBeYGX02WVpPYAyv0
38UFjXQpQBG8oKXHxDlZLB5kV6a7V4erPXd7KIytC5G1HAl34B0Yg4MxIYuYf2C3yPHFM1awKsoe
JeuCOXNym9EDZZFvNnUtALHrK6KV1i153dU5CB43gXNUDklJmnEyU8gWw18Ap9LJYI2NPv38C0eu
eW3D6S2D6Q5LtvmrEQjIGApdZHD+qyMN5tYZbShXTCXtrTdIIwzFNZSA8Vu8wTbfGI9xuEkXuqL7
gywZHsui+GYDQdaOsCNrvLXg7ER5v6HS4iUYtBum8bM/SD3G8ZlXd9J4/Qg6L6d4Hw66T4AUc4KO
BTqM0dpXZV4sjzJFvTu6/47m+LdmPQrgR5aCPr2ZDBSjAOG0skDINJ1Pmh9a4A9USfqfUpu9SCaQ
silJP2t1yBfhNVT0wJOWLJVVH/gzxZpeU0rrujYgPnGRCVGp6bH9MPYHnbZ0pX0kPSqwaWRg/PR6
kETI0isNGZIaO9rnbN1sqjFJn4LAYdl2lURyx70L4YLM6EKsjwsRZES06sD7JOrjtHZUiIigIllw
1ZHQ2EYjIeiLqJcgbZkKnNj5Um9tt2DPPIraSkLcI4pe0wUXg3UxQYvZ63TU/VyV
`protect end_protected
