-------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 2.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard
--  /   /         Filename : gtwizard_0_multi_gt.vhd
-- /___/   /\     
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module gtwizard_0_multi_gt (a Multi GT Wrapper)
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;


--***************************** Entity Declaration ****************************

entity gtwizard_0_multi_gt is
generic
(
    -- Simulation attributes
    WRAPPER_SIM_GTRESET_SPEEDUP    : string   := "FALSE" -- Set to "true" to speed up sim reset
);
port
(
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y0)
    --____________________________CHANNEL PORTS________________________________
    GT0_DRP_BUSY_OUT                        : out  std_logic; 
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt0_drpclk_in                           : in   std_logic;
    gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt0_drpen_in                            : in   std_logic;
    gt0_drprdy_out                          : out  std_logic;
    gt0_drpwe_in                            : in   std_logic;
    ----------------------------- PCI Express Ports ----------------------------
    gt0_rxrate_in                           : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    gt0_rxcdrlock_out                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(19 downto 0);
    gt0_rxusrclk_in                         : in   std_logic;
    gt0_rxusrclk2_in                        : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gtprxn_in                           : in   std_logic;
    gt0_gtprxp_in                           : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt0_rxlpmhfhold_in                      : in   std_logic;
    gt0_rxlpmlfhold_in                      : in   std_logic;
    ------------ Receive Ports - RX Fabric ClocK Output Control Ports ----------
    gt0_rxratedone_out                      : out  std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    gt0_rxpcsreset_in                       : in   std_logic;
    gt0_rxpmareset_in                       : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    gt0_txpostcursor_in                     : in   std_logic_vector(4 downto 0);
    gt0_txprecursor_in                      : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt0_txdata_in                           : in   std_logic_vector(19 downto 0);
    gt0_txusrclk_in                         : in   std_logic;
    gt0_txusrclk2_in                        : in   std_logic;
    --------------------- Transmit Ports - PCI Express Ports -------------------
    gt0_txrate_in                           : in   std_logic_vector(2 downto 0);
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt0_gtptxn_out                          : out  std_logic;
    gt0_gtptxp_out                          : out  std_logic;
    gt0_txdiffctrl_in                       : in   std_logic_vector(3 downto 0);
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclk_out                        : out  std_logic;
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    gt0_txratedone_out                      : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txpcsreset_in                       : in   std_logic;
    gt0_txpmareset_in                       : in   std_logic;
    gt0_txresetdone_out                     : out  std_logic;
    ---TXPI---
    gt0_txppmstepsize_in                    : in   std_logic_vector(4 downto 0);


    --____________________________COMMON PORTS________________________________
    ------------- Common Block  - Dynamic Reconfiguration Port (DRP) -----------
    gt0_drpaddr_common_in                   : in   std_logic_vector(7 downto 0);
    gt0_drpclk_common_in                    : in   std_logic;
    gt0_drpdi_common_in                     : in   std_logic_vector(15 downto 0);
    gt0_drpdo_common_out                    : out  std_logic_vector(15 downto 0);
    gt0_drpen_common_in                     : in   std_logic;
    gt0_drprdy_common_out                   : out  std_logic;
    gt0_drpwe_common_in                     : in   std_logic;
    ----------------- Common Block - GTPE2_COMMON Clocking Ports ---------------
    gt0_gtrefclk0_in                        : in   std_logic;
    -------------------------- Common Block - PLL Ports ------------------------
    gt0_pll0lock_out                        : out  std_logic;
    gt0_pll0lockdetclk_in                   : in   std_logic;
    gt0_pll0refclklost_out                  : out  std_logic;
    gt0_pll0reset_in                        : in   std_logic


);


end gtwizard_0_multi_gt;
    
architecture RTL of gtwizard_0_multi_gt is

    attribute CORE_GENERATION_INFO : string;
    attribute CORE_GENERATION_INFO of RTL : architecture is "gtwizard_0_multi_gt,gtwizard_v2_6,{protocol_file=Start_from_scratch}";


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

--***************************** Signal Declarations *****************************

    -- ground and tied_to_vcc_i signals
signal   tied_to_ground_i       :   std_logic;
signal   tied_to_ground_vec_i   :   std_logic_vector(63 downto 0);
signal   tied_to_vcc_i          :   std_logic;
signal   gt0_pll0outclk_i       :   std_logic;
signal   gt0_pll0outrefclk_i    :   std_logic;
signal   gt0_pll1outclk_i       :   std_logic;
signal   gt0_pll1outrefclk_i    :   std_logic;

signal   gt0_mgtrefclktx_i      :   std_logic_vector(1 downto 0);
signal   gt0_mgtrefclkrx_i      :   std_logic_vector(1 downto 0);
 

signal   gt0_pll0clk_i          :   std_logic;
signal   gt0_pll0refclk_i       :   std_logic;
signal   gt0_pll1clk_i          :   std_logic;
signal   gt0_pll1refclk_i       :   std_logic;
signal   gt0_rst_i              :   std_logic;
      



--*************************** Component Declarations **************************
component gtwizard_0_GT
generic
(
    -- Simulation attributes
    GT_SIM_GTRESET_SPEEDUP    : string := "FALSE";
    TXSYNC_OVRD_IN            : bit    := '0';
    TXSYNC_MULTILANE_IN       : bit    := '0'     
);
port 
(   
    RST_IN                                  : in   std_logic;
    DRP_BUSY_OUT                            : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    drpaddr_in                              : in   std_logic_vector(8 downto 0);
    drpclk_in                               : in   std_logic;
    drpdi_in                                : in   std_logic_vector(15 downto 0);
    drpdo_out                               : out  std_logic_vector(15 downto 0);
    drpen_in                                : in   std_logic;
    drprdy_out                              : out  std_logic;
    drpwe_in                                : in   std_logic;
    ------------------------ GTPE2_CHANNEL Clocking Ports ----------------------
    pll0clk_in                              : in   std_logic;
    pll0refclk_in                           : in   std_logic;
    pll1clk_in                              : in   std_logic;
    pll1refclk_in                           : in   std_logic;
    ----------------------------- PCI Express Ports ----------------------------
    rxrate_in                               : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    rxuserrdy_in                            : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    eyescandataerror_out                    : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    rxcdrlock_out                           : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    rxdata_out                              : out  std_logic_vector(19 downto 0);
    rxusrclk_in                             : in   std_logic;
    rxusrclk2_in                            : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gtprxn_in                               : in   std_logic;
    gtprxp_in                               : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    rxlpmhfhold_in                          : in   std_logic;
    rxlpmlfhold_in                          : in   std_logic;
    ------------ Receive Ports - RX Fabric ClocK Output Control Ports ----------
    rxratedone_out                          : out  std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    rxoutclk_out                            : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gtrxreset_in                            : in   std_logic;
    rxpcsreset_in                           : in   std_logic;
    rxpmareset_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    rxresetdone_out                         : out  std_logic;
    ------------------------ TX Configurable Driver Ports ----------------------
    txpostcursor_in                         : in   std_logic_vector(4 downto 0);
    txprecursor_in                          : in   std_logic_vector(4 downto 0);
    --------------------- TX Initialization and Reset Ports --------------------
    gttxreset_in                            : in   std_logic;
    txuserrdy_in                            : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    txdata_in                               : in   std_logic_vector(19 downto 0);
    txusrclk_in                             : in   std_logic;
    txusrclk2_in                            : in   std_logic;
    --------------------- Transmit Ports - PCI Express Ports -------------------
    txrate_in                               : in   std_logic_vector(2 downto 0);
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gtptxn_out                              : out  std_logic;
    gtptxp_out                              : out  std_logic;
    txdiffctrl_in                           : in   std_logic_vector(3 downto 0);
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    txoutclk_out                            : out  std_logic;
    txoutclkfabric_out                      : out  std_logic;
    txoutclkpcs_out                         : out  std_logic;
    txratedone_out                          : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    txpcsreset_in                           : in   std_logic;
    txpmareset_in                           : in   std_logic;
    txresetdone_out                         : out  std_logic;
    ---TXPI---
    txppmstepsize_in                        : in   std_logic_vector(4 downto 0)


);
end component;


    constant PLL0_FBDIV_IN      :   integer := 4;
    constant PLL1_FBDIV_IN      :   integer := 1;
    constant PLL0_FBDIV_45_IN   :   integer := 5;
    constant PLL1_FBDIV_45_IN   :   integer := 4;
    constant PLL0_REFCLK_DIV_IN :   integer := 1;
    constant PLL1_REFCLK_DIV_IN :   integer := 1;

--********************************* Main Body of Code**************************

begin                       

    tied_to_ground_i                    <= '0';
    tied_to_ground_vec_i(63 downto 0)   <= (others => '0');
    tied_to_vcc_i                       <= '1';
    gt0_pll0clk_i    <= gt0_pll0outclk_i;  
    gt0_pll0refclk_i <= gt0_pll0outrefclk_i; 
    gt0_pll1clk_i    <= gt0_pll1outclk_i;  
    gt0_pll1refclk_i <= gt0_pll1outrefclk_i; 
    gt0_rst_i        <= GT0_PLL0RESET_IN;
      
   
    --------------------------- GT Instances  -------------------------------   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y0)
gt0_gtwizard_0_i : gtwizard_0_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RST_IN                          =>      gt0_rst_i,
        DRP_BUSY_OUT                    =>      GT0_DRP_BUSY_OUT,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt0_drpaddr_in,
        drpclk_in                       =>      gt0_drpclk_in,
        drpdi_in                        =>      gt0_drpdi_in,
        drpdo_out                       =>      gt0_drpdo_out,
        drpen_in                        =>      gt0_drpen_in,
        drprdy_out                      =>      gt0_drprdy_out,
        drpwe_in                        =>      gt0_drpwe_in,
        ------------------------ GTPE2_CHANNEL Clocking Ports ----------------------
        pll0clk_in                      =>      gt0_pll0clk_i,
        pll0refclk_in                   =>      gt0_pll0refclk_i,
        pll1clk_in                      =>      gt0_pll1clk_i,
        pll1refclk_in                   =>      gt0_pll1refclk_i,
        ----------------------------- PCI Express Ports ----------------------------
        rxrate_in                       =>      gt0_rxrate_in,
        --------------------- RX Initialization and Reset Ports --------------------
        rxuserrdy_in                    =>      gt0_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt0_eyescandataerror_out,
        ------------------------- Receive Ports - CDR Ports ------------------------
        rxcdrlock_out                   =>      gt0_rxcdrlock_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxdata_out                      =>      gt0_rxdata_out,
        rxusrclk_in                     =>      gt0_rxusrclk_in,
        rxusrclk2_in                    =>      gt0_rxusrclk2_in,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gtprxn_in                       =>      gt0_gtprxn_in,
        gtprxp_in                       =>      gt0_gtprxp_in,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        rxlpmhfhold_in                  =>      gt0_rxlpmhfhold_in,
        rxlpmlfhold_in                  =>      gt0_rxlpmlfhold_in,
        ------------ Receive Ports - RX Fabric ClocK Output Control Ports ----------
        rxratedone_out                  =>      gt0_rxratedone_out,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt0_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt0_gtrxreset_in,
        rxpcsreset_in                   =>      gt0_rxpcsreset_in,
        rxpmareset_in                   =>      gt0_rxpmareset_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt0_rxresetdone_out,
        ------------------------ TX Configurable Driver Ports ----------------------
        txpostcursor_in                 =>      gt0_txpostcursor_in,
        txprecursor_in                  =>      gt0_txprecursor_in,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt0_gttxreset_in,
        txuserrdy_in                    =>      gt0_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txdata_in                       =>      gt0_txdata_in,
        txusrclk_in                     =>      gt0_txusrclk_in,
        txusrclk2_in                    =>      gt0_txusrclk2_in,
        --------------------- Transmit Ports - PCI Express Ports -------------------
        txrate_in                       =>      gt0_txrate_in,
        --------------- Transmit Ports - TX Configurable Driver Ports --------------
        gtptxn_out                      =>      gt0_gtptxn_out,
        gtptxp_out                      =>      gt0_gtptxp_out,
        txdiffctrl_in                   =>      gt0_txdiffctrl_in,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt0_txoutclk_out,
        txoutclkfabric_out              =>      gt0_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt0_txoutclkpcs_out,
        txratedone_out                  =>      gt0_txratedone_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txpcsreset_in                   =>      gt0_txpcsreset_in,
        txpmareset_in                   =>      gt0_txpmareset_in,
        txresetdone_out                 =>      gt0_txresetdone_out,
        ---TXPI---
        txppmstepsize_in                =>      gt0_txppmstepsize_in
    );


    --_________________________________________________________________________
    --_________________________________________________________________________
    --_________________________GTPE2_COMMON____________________________________

    gtpe2_common_0_i : GTPE2_COMMON
    generic map
    (
        -- Simulation attributes
        SIM_RESET_SPEEDUP    => WRAPPER_SIM_GTRESET_SPEEDUP,
        SIM_PLL0REFCLK_SEL   => ("001"),
        SIM_PLL1REFCLK_SEL   => ("001"),
        SIM_VERSION          => ("1.0"),

        PLL0_FBDIV           => PLL0_FBDIV_IN     ,
        PLL0_FBDIV_45        => PLL0_FBDIV_45_IN  ,
        PLL0_REFCLK_DIV      => PLL0_REFCLK_DIV_IN,
        PLL1_FBDIV           => PLL1_FBDIV_IN     ,
        PLL1_FBDIV_45        => PLL1_FBDIV_45_IN  ,
        PLL1_REFCLK_DIV      => PLL1_REFCLK_DIV_IN,            

       ------------------COMMON BLOCK Attributes---------------
        BIAS_CFG                                =>     (x"0000000000050001"),
        COMMON_CFG                              =>     (x"00000000"),

       ----------------------------PLL Attributes----------------------------
        PLL0_CFG                                =>     (x"01F03DC"),
        PLL0_DMON_CFG                           =>     ('0'),
        PLL0_INIT_CFG                           =>     (x"00001E"),
        PLL0_LOCK_CFG                           =>     (x"1E8"),
        PLL1_CFG                                =>     (x"01F03DC"),
        PLL1_DMON_CFG                           =>     ('0'),
        PLL1_INIT_CFG                           =>     (x"00001E"),
        PLL1_LOCK_CFG                           =>     (x"1E8"),
        PLL_CLKOUT_CFG                          =>     (x"00"),

       ----------------------------Reserved Attributes----------------------------
        RSVD_ATTR0                              =>     (x"0000"),
        RSVD_ATTR1                              =>     (x"0000")

        
    )
    port map
    (
	     DMONITOROUT             => open,	
        ------------- Common Block  - Dynamic Reconfiguration Port (DRP) -----------
        DRPADDR                         =>      gt0_drpaddr_common_in,
        DRPCLK                          =>      gt0_drpclk_common_in,
        DRPDI                           =>      gt0_drpdi_common_in,
        DRPDO                           =>      gt0_drpdo_common_out,
        DRPEN                           =>      gt0_drpen_common_in,
        DRPRDY                          =>      gt0_drprdy_common_out,
        DRPWE                           =>      gt0_drpwe_common_in,
        ----------------- Common Block - GTPE2_COMMON Clocking Ports ---------------
        GTEASTREFCLK0                   =>      tied_to_ground_i,
        GTEASTREFCLK1                   =>      tied_to_ground_i,
        GTGREFCLK1                      =>      tied_to_ground_i,
        GTREFCLK0                       =>      gt0_gtrefclk0_in,
        GTREFCLK1                       =>      tied_to_ground_i,
        GTWESTREFCLK0                   =>      tied_to_ground_i,
        GTWESTREFCLK1                   =>      tied_to_ground_i,
        PLL0OUTCLK                      =>      gt0_pll0outclk_i,
        PLL0OUTREFCLK                   =>      gt0_pll0outrefclk_i,
        PLL1OUTCLK                      =>      gt0_pll1outclk_i,
        PLL1OUTREFCLK                   =>      gt0_pll1outrefclk_i,
        -------------------------- Common Block - PLL Ports ------------------------
        PLL0FBCLKLOST                   =>      open,
        PLL0LOCK                        =>      gt0_pll0lock_out,
        PLL0LOCKDETCLK                  =>      gt0_pll0lockdetclk_in,
        PLL0LOCKEN                      =>      tied_to_vcc_i,
        PLL0PD                          =>      tied_to_ground_i,
        PLL0REFCLKLOST                  =>      gt0_pll0refclklost_out,
        PLL0REFCLKSEL                   =>      "001",
        PLL0RESET                       =>      gt0_pll0reset_in,
        PLL1FBCLKLOST                   =>      open,
        PLL1LOCK                        =>      open,
        PLL1LOCKDETCLK                  =>      tied_to_ground_i,
        PLL1LOCKEN                      =>      tied_to_vcc_i,
        PLL1PD                          =>      '1',
        PLL1REFCLKLOST                  =>      open,
        PLL1REFCLKSEL                   =>      "001",
        PLL1RESET                       =>      tied_to_ground_i,
        ---------------------------- Common Block - Ports --------------------------
        BGRCALOVRDENB                   =>      tied_to_vcc_i,
        GTGREFCLK0                      =>      tied_to_ground_i,
        PLLRSVD1                        =>      "0000000000000000",
        PLLRSVD2                        =>      "00000",
        REFCLKOUTMONITOR0               =>      open,
        REFCLKOUTMONITOR1               =>      open,
        ------------------------ Common Block - RX AFE Ports -----------------------
        PMARSVDOUT                      =>      open,
        --------------------------------- QPLL Ports -------------------------------
        BGBYPASSB                       =>      tied_to_vcc_i,
        BGMONITORENB                    =>      tied_to_vcc_i,
        BGPDB                           =>      tied_to_vcc_i,
        BGRCALOVRD                      =>      "00000",
        PMARSVD                         =>      "00000000",
        RCALENB                         =>      tied_to_vcc_i

    );

end RTL;     
