`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IGOUWam3utmfnHmSGpINKp1TTk1PWR1CXkvtcqb4kTkTUgGwxq7FbZqSBxxGUeeRYzzIBvOk5pMM
ngzo7VIIU3RcVfOS8oYSTezf483Tt0IQtK+MS2dYHA5q30qwV6KgufZ3dgFklmZA3LNVU/59/kuC
VjyvMLqFeh4dP9OD2pmdoL+nP/AEh6KPQlA3qV51AsLz/CdtkDaTPWyl7fXQ+KpmKDb4vMmI4eln
dHAisbbD7idDi9kAnylncb/elFoXT+UaVDwJDk6u1ZTChdH1O2rPdL8eFK2tvGS4c1aSUzDKHAOO
nxr8aG8QMAC0/Um+D+WumXmTwVsU6U6pRrLapg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
E8Eg4M4oHZ6ttL2oO83cjIjRvxKoYRs7rQIOKt8Eu/AMqZIpCyh/dpBXqSr9UsbswBtDUcPuQWmY
fEmahfWPYMwEPL4Rbl3Sl0hEJkkdmRl5FZohwiGgkTJMZmkmggN44cak1eP71Xj8r76i8wpxxF4P
P+3D+qBsHU30qWYIJn8=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
czCO8K4kQRIx6BQKyGIoOxiSexcyCBYhcvhvPUHcUbEC3XyArPWosTrmFn2iPrEa3c0QY1gxh6ES
xK89hdSKmHgDFs4GEVJLjcP8R3Jsm1cjfjae3RxJwD1wbeQSbJ8JqjazK3zQrveGg0ngQpghqF2i
wqS2MiY+jN64ITi8L/w=

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15040)
`protect data_block
VwSfIV/TCQiKhUu1MkKled+CARVt3v68xiifNN1VpGGRuoYGg7KiPXWgK7GwIPaNxdmUmXkirRA5
6Toz79Tq3KK3aX5YMYT+c0vSa0FdIsWvg2bvfCpV8Ugq0KWkrq3mhl2FkSr2y99TCEgWMwjkvQnP
sdBbk3CNAojT+AfOd9Vw8wjF01NWNQPeyS+WUIOH2DLTnrONqUjqPteTRJ+qOgTOJJ4eL+G11mX4
4ZdRtutHV9v7u5eVYUuGp6jjjU47SsTT0blqNQPckqCNWtP+qXn9r4PiRffmtkRaLQ4QQ39zlHzr
iZB8OVZPDCXoPd/DQ52XEC7P2SmiQkjuPh10tD/9JV5ZRQcpw6HowVm1rK4wEjgkfia/zHyIRFUg
ZJF2PPe3jMGst7xLKq4XW09phVGVO7e7fw/hcbmiq7xV4vcDg8lSDEbqh5G9kLNnDbUK0yaGSh2N
ciDYkf+M4S+adR9UWxASZmWnaznDjMi7ZSOpOLYOW72qIIUXl1y3bqyQIvK2RXdpmk9QRWTAONOb
8BpMoSkOYkTx15O8btvb0P0AQ9kAsUPxCBewDb6asEbhNs7sCdrSL8FIuvOW8G7+HCv0D86ZZwck
5d6ZUBa4+kX1ENC8zZwCTS3k68LMRifrPQ0cRspAJP5IFbvdeh5dRPM+9H+GC2BNqjA3ElVa1DQ6
3Uwy8zOxuBExiYmG90wDnwCa7TWPpqHSyhyioOHK8y4aNjlqK8RmVZv0AfiqKIp5OscKpwojD7IR
BlvGtU8N7HlaUN7R5rJ06lj/kjPJ2WOGPsc5BK0TCOA2utv+UEWrQMSUfF0JhIT4Qz1DQB56FEza
CD8a4cSN8SgEY91wQqusda+zZ+tEgI2jK7aBfmaI2ypgl0qusMLAr022zun+g1kCN/6boL3fUEUo
wucN7ykLG0Wz+68Afbd9ziF3bgyfxMNTtJMGs1PSaVy1CNtJBUjd2eVeYdz9HfIMkX4ws9VOxmx3
0ChoTz7xL2jgy/2UQzlnnbAJTMCsbhpcVtK6x9WXibjs0WJHmr1mA3GA2zVqUak2Sliq+N8DZgL7
WayV6ap3A0Mrssl/tkOx/1midjL/wN1UfQ2+SfFlpvseUHGhhHHp4sK57oe9E3ZxuNEMQ7Hs9RS9
qqVbnWz+hYrte5BpDhtVsUPVPosMSPT5tKv0ktyIMFimjj+N8sXzTyrIbBt8z0xFay1HzLy85m+5
bsQ3tqPOyA0q8kf0a3kNPhi3KkQuI2JZg56wWo9XhGMNslmStAttPvhzBSqXh4qu9pP+TspPCDxL
oNh3EEUVLWS+1aH+tfSEUNWzk7uasckRXq8K9z7QGcgWGAnKk2gFukQyuKjMgoo+UwbkC2SwSTVy
iZn+soXLMxT2pdKkBttzewJJZIa4opqoSCL5lOASa15ZMYhiHldUij+/Dj7Oo1g0UPQv6peLiDjQ
K/lBaUW87dOfJC9Y9qer2C1s8EcME8WywV77h2xP5frmpdbuxUTX79TtAfLh+1+dmmxdHFGCSC0j
BQlIy5ghbDqYTgyqISKGHsrj98/lWS0+UyHDSvsBB+p7x1WQuXc5JGIxVjJCl3iUI9hu4ik6p/qg
ahG4Bpap4VCHeNv6qqJF/iINEElgSlKvqwyGKoMe1WjpISrtrMUD8TN13GuYm5+uOcTqUdmmc2K0
0fCoIL08b63gBpNuIdlJHX99b1jfaLsqljoPrL4UcCHB5X5VURTs5015mBr3KQKPoCVVwq4ZzPUn
uGeptNS2FFrJ+GCQkyoupa/LsU2sg80eEcg4Z4pCzwRWBkbpyi/B86jYl6gPXjUvdl0gyAHliLRw
n9L7RA49csl7JvZzdUvjPBJKMKPp11Jk1jouQ6qs3moUfdBS1EsC9ryW6yxcKae6Dp/oRxqVHUUT
iF4t57cRoZS/vln1VXSIv8Hslz78IL9V44JGk7ZarpSwjiHDtSKa0aeLFBT49M527cL4jTw55RKH
KMuJ58edGAmf2FbZDESgv5G93muQCjhzpzcEy+JV8fj8yYjt5WnVmwT9hzsMHNbpGrJf0JMpmQJi
2gAf4DQOzS+a7n9yl7wpWYjFwhkb7E8MgijjFuYKpEaEC+YcyGFjxcOXpsyEuw2Fwf5o/X9xaKdD
YxxY+he/21GAQDUWcs6LXasro0MhrKjkVVrAb68qF+uDVWi1xxqRetFjdk2unbVPZQcMzZVN5rY7
KznCQTmJIy1/YF914QGl4tQGHzcoJf07g4kL/OryEh0UmXYmKey4VE6mDcqzu36cP1FbynPQrYEh
aatxW4iI+uByUwkKs0ZGkLuwqUYEN54UDVZsZW2F23O2a/NHyD89gXhTMEs7X4A0snRTxC0fvHGf
UYfgG6WNdNnnESbaNvoXbTztirYGUOUNTml0DCK+K9SXpa6XtZgLE/P1pcZQORGKUpFTaYb4do5r
z1i2hRjgzVC0k1LcElsRe5ww6XiZfB9tuzMoY6PNkO8liyO5pEGGi2adgesZediSYNLa3xEKwakC
BLOtgpUPTXNefdkKTdhYomMx2ShIwn0aNVH2p5niuN3/V2+zhD+z0HiYlEGo2omKOfdagAAR1kOj
ds8r4FkqAPR5dp4xT6Z+MpWd+q+dDjurpdfB52fq5qsg6FpmE88ErB4EtcQgMGozgj3qUSmMaMyF
X0G9SYfo0kWk14akaonFteuyY0l3FAvAenaUEpasot5jbjT/4WXNRLjLqQ4rhpwpHabew7zbj0JI
Rhd21u6X9yqp7i85TD2eyxOpsikiJCVbEErhAVosx+CUOS9fxmuS3DdkQLxbntOo9MP5+xPuHvlo
KeZJhMFwhkFoZKRjniq2MNGXd3mqHnZ2M9N8QYOPdAgz4AWiZW6sQiIUR84wikFnWD6/2ZHq9knA
IVGy20FB+L6Zplz6P6lg9MT8LuFPUD2ZUvChS5f+BOvhSRrmoZZ2FTC7adWPjMNuuR12o8CbqVXt
lMJTyXgc5GxftZ3dgrc/0TFdp4sqnodFmXIjdWyoV5Tm3CNxR/s/ZUEJr3P0Da7g9NCMHfSovKV3
w6IS/lmUcC1EplZ+i3/j6ZTT3G8F3wqgHd5PBYwNZUv6yEOmkoAasZIK9SVyyMEBJS7qipscpntZ
jn/IRP098JxesSDLtd4k8F505NLaQiLk/0S1xZ+gEtreN7EicJ26CMH1xwHCHjmu/PXSYE5JP+ZR
PuP1FL4drktdDFpx+Pd1hekgFgBPWbTRehT2R4GoKcAXN6LL0BfJWSIeSZF5czGwILm+sN+W7i0T
j8eynXxh97fW5/MCTD1W5dvAVC+fcaEo0bLV5mKtgC1SGrKSi0iPGA42iK2wpP3YnNpYp0uWlBch
XOfc1bm1jgF859I3C5rd3HUYxf47Hf3+Gfd2SwYtNq+rfPK1BEU7lLofBn7LdQg87FIZ+3nvPgr7
xxUARpepRtH15uJOk68qLLzUF58UsB4VlV7/a8Z8nFK2PHESGmJjn3ifrKjg6cdXH72kMas0HYdV
kp/QW4vRGWw3U3v5sE0zIoRkWbQ53ZTk/NZXgDnDzXxAk9wHLLHVA/AOv7ime3SiWdzahBXmqkUR
+o1LOWSZx5fu5Z9lyNuN41T7gsSybPWxBnD5gygq0f4XUfrsiJH5YYuixef/jmswVbqeteCkyvlc
Q0jkiHIDxT68DI8+ulTJCqdKdYd7ZkuphuAeSml6GlOb/g2vfSaPjebnLXdQ8v8qTuCt7b9iWrKA
D46Ix+Pn4QB8sPTZ4W3PvEiaCR0to+YRp93r48iqr6Rmt7MzdwGPWs1bJgtCeuFrZzm/MPsuc9Zn
T6AXdacfzubwn6xryhRKe/mOJUjUdhbm+O1ZJRZ3EJxJw88/7dpVeiAnxFWeSSSbL154fnEJ3wsJ
McNsbI2wxdS+JMtjU5UpudPs/CyMFCIjVdn6lb1Z7UbUay5BGq1WFSr3AtCQ/0CAqlII03KA2sVm
ilNmBeQl2ENB1LuJSM9GF6RyW01RiNcELo6sMclieRYt694PLX6CmJxv94GGAMCYr+e/FUZVXS/L
YWY7c2nCPyVdy6I0IvDi0r0oI2UfXXHhryvKIxUMAJjg1genLdywEHgi+Q5pe2q8PnNpQm3SX3r9
m4XwWHL+cj9ndBMkU9BrI9oWT08wlcp8nMVv0FgMJceO3HLy7ujcYwYUu1gbCyKYf4mffpTvWU9a
26yLncK7hvnJqynz3lRllUyD5MKQwJ5C+9+W7hhwbi4cqY59XGKmhyDgaYUe5HH6kO5mB75ernLa
tAScJOq/Ba+8XqDsel1srsNaaSTwMD4VuZ+M19qEXtrMHjMKyc6OSrMZJaJe1qd/D0KxU9uP0GDf
fUmvrWj572Qq/OKUm9xPbXyS7f7KFNiY4tPobkESEJZm1/pfuFEkR6ifAODN4MwXs1wpHoG673ks
Hfc8236+GzNOcZMnRSNFrOs8azdGzvmZvIwr1htlbOv/w32KH8/Nhb5WH3IxjzldypFPP1euuKSq
E332NB/60T+R7zpPXASBToBFnUmFodoXLmcXAffT3gSsVhu4F7nzJTBCh+dLo2wWNZpg8L5sI/Bi
CEkacJNTrmgrubvZ25O4f6TTLxbcaWOCFOa+YtjT15Qb1JdT1/RX7DJV2rfMJLH3Hm68u1F7fhra
E0cIeeUA5ZxcHzwIlaabDL+KSUg3ZCWoytffrzBF+P5e1jwvvds/5tvsk+YeolIjjIfRD5tNxHwJ
mYNzg9A8FuweXneqg+4WFP1vNogTSU7JekpsWVZSiBMmL0FxNjqNHLI/V9LgMNXpH9cjOIRwMn1c
MVHaplzAznXLRhWnKBOufGUZvaCb5Vg/Fpgrfy3Y1YBDMV365qdxXkFnMhQLT1nfUD0zmqH1f5iE
5b3QrsbPg/Il22eFFAoh1KN2232dL9eGPPtUaMOIG/73Ifq9vHMtHUT/VFr4CwoSvMybSQVx6SOb
TbpyBUl8QO6l36s84NNXOAJzM4+DP3EbXuYcBJ+IUEWhqkkotku7MYH+cgrpFrGpPIEQtYXoTRFt
fUSm05wGwtixSlEyr547h2ODuEJlircN9trluidUi1EKFGJx8W73x2OrlBbnMfvp/ATLyCNanE3u
vCf9ft/+Op88bJPu90YFev3TDPmeS2+pw8yrGslhew77I1vmVUFCdkxDZLIJUNB3vK3HXFUiVAyq
d0jmdhOpTV4Mzfq0Yk56zl6MXD1fnmXi+I4HCIu1UMSu5nAVRA6Bv91GhUsxXqN3a+P9DrtObXHj
cWHAy2/u0X3BqUO+CQgjIrLSsAqItlTTAfwOP2+MtbquTF3xmBM2ww+FYBdDoDBDLeBxHAE0M+n+
cNGp0RbDhp04Vyxkk0x+lx7ym/1rhk11f0nSpxH5ctyWRikECbKm9tvwPjnfhYD4z4M6gd0OHwbl
1PoyMdnVFD/BPXuOsvirLODaR1laVNfQWPLIYikhkc2FkRMXZYB4IGE0Xp3KzU8EYrjVvfCHesNA
FNl8iC0QJ09M0cIU16GwndU/c4rNh2gJgF7ie8V6jYLvaiVlMxZDkEj/9sPvbnpj8Z3qdPYbOag9
y8/W67MtzmvkHJiAWu6Do7jKtgMVuvZoV0Ht2QpkpzNb73ezAydG/T8w1tXl8MN2dTolP3wZX7Jd
+S98ts/31grnMDz1jn2NuJhMbZI0B0j/9idqWVpcstzlZO77mN3l4GCTHShnCfJ7f33oWYPiPyJ2
YCgm77EBaSpUdyBJcvSBuIbluv00p7uUv/RkNhc9ZgOb3Omoe752Xx6Aq3XH2oqXPNNwCDTpCXEL
xi/Ds6hp1T7DoOASzSNP3SwrA7aqMQzOWsgAmRmUaZ6xer7TmqbsLTBF4fFON5FWiJsiSDztrbrN
orR2YHVpnKRB1DVGyBvVEJPu+pC9eVLEAXPqJqtGeh1AJZOAFHoDLxM5auYyPvx3R6quusERIYjs
uaP298EsU38qoD8rBKdritxsJ/bmp63BWOEPBJmD3Q0gOLI3r9XocjEbjpPQpdWXqg6awX6TqLAR
q8aP0Z4Hr6K1RiD9z+SxNEz5wPkXmDiNH9z4vt9JhlYxPisuofyjcSPL1hdVmNccGnSvEBJ6nYoW
hRuzthCA4nUld0gF0JPpAbXqNNDojFJBZqy0gQ0/6JyWqWmF/EoxJjxkkOgqZRT0rmW5qpZ3B/Uv
llpwo9Xa61T2tlET0CB6mg5AIiXTxV4IP417NYYFk2A2Hum9kjscYJBr4ZtkLGN0lDo8R8gXpsG2
D0zqBkI4wJmRR+UgXwy3tYUXkj02gN3HSN3Oid3kGvwSlGm2zmWi1EiG4IMG5PncCpkp87wgKgsd
SQYOXGgG4GlcaJkXyc16QovmQXjHCzPEFYOqhHhLxqc//fDuUH4XZLlIjg0lxbAYbDDaw0uZ7gMC
MJvzaqrthH190/cVASKg8qdHSIPomKoJkWDLQ95MCRIk49RUZepCiKTPrZZAZXnHZtl7GH6LSuSO
q09N+x2ixvnGQx/qU1HRH0BpTrN12HXYq3QZIIWG8tV9rGICGbuQiO+h5O6CFIFq+b/W6K6ab/RU
3S6qkHpcid8lZXt6j9gZt30O9BIdVn0TcHErbjHogMN/M2d+SLsy3Lx6MeT7DCZbX1g0wV2O9onp
oA5pGVgGVicZBzUJhK21oBqRMbvKyTDsrLnaVy/vvTGKOAWumHMxV6PCPLQYzoemFWxvSQMhvlb8
Pd/yptu74TP6mkAfz/mUpR6LxGRxOgx/9owpVh+UHEuAmbxhH2kYQHhbCNGMPmrpleyACyn/nvhe
tW/ZS3zS1ul2w9pD0EgSBz70+QDLhAlQCLMaaew1XAqZ9SnfP5W1krTjCJL4Ud81/Y+e1wtBugUB
04ZU2oXTXyZy79AvZDoB9HEsWTJ0GI7EZ1DtshACCno2hBxg8TLtDQrfsiHgZUXwyR6fF5GC9KDM
93U3dMaBTJLMszUHzO9t7IpBDDGRX3qm/Z/HbdBj3q+cGYu0K47iODeeA1InJoBKqUQRZBSd82S5
HnmnMpEH/bCKuagOWtm3hPx3W4OYhwulE3rbhiBE6qDKldq2UHyttOlnSblbUBQW3krnMSfz/z5X
2Lm/G4hrcqNWQ55KbWW7ai6XR/xhLWQoqDZVl9BUV315oZJQ/VzOIBH+ueZOH6WhcbZF0OUvqX5F
5R5sW6IMHIxDuJ8+36POL3qdUCNRGt93wf2q7KMYOCI6U6+5x1V3SGbaDO3cdXq3npNIBoUzUEV0
tQRxp/cT3zNpj1sHM5s4PL+QKoYdK63bTKHLkJwEXLPslTkZIEVQUsK71ureo99HYUvqjMVDu4Bl
EajwY2ySmlSoz1OIGbuhcS5pq1waxgk/3sYj8/uH4c0ATLPAgiyerbVQASzdlaCROIV8r92IKSvw
InEDaZS9O+qYjYfoxohR4Y4ogga8NbaI9BYO9sTUyKDspaY1tVJsU+Wd+JpuR2G4GteoYd0LtVjb
9vRzRXvCb1r6Y6yZu4CVgm3zQtPe6u0+qkrm27h34+yIw9lSGUBHAAnHyQJRHb/CPd4Ihyuj+aBR
G8otcmfllJE4kwHTv4sqFhbqHzFAC8D5hxr32nqJxWsbimbHvV2K4wYg9dtIUmq8CND7sP4MNv9h
4d78oIjMICMIrP5r/6clAFrYyaoDIKN9LnLxwfuhd/SjVHOqOHNx9k1sDayezNCKPDnIwloM7FUq
o2vK+GOvOFNj1i9zjyuPvqzakbVwFEcjXkLbG+o9hIn5uBnkKHbG5+VbevhqA57UL9rBPsMa1Ztm
e8NwRKI0QX5zSDy2nuFpRxnai7cfG5bojdv7fxpwrRrpFwK2jdFSMAviR/IHtZk/HDiQOmA5GSPT
kh+VhqQd5qsDWGLN71/6tHUk5P99F8jp49uKoac40eNVPYGKIiwc0yRX6J6wEpysbg3utl2PpG9d
nNWsuLtNuir8YX/xxP85WPZgfVc6cjm8b873xXCNYSGVi85K3lgnB5kqPpyzyWJmLCt1kSvGzA30
ddL++qSN4Kaym1fs1z7pmalreyuigW3Rk37ZGng7kkDFrDTElO9vL5ROsg6TnHFMgN58+HK6I8Iw
ESoTDGNPD7xnKd9XhraVwpQn1slCxDHiNuEHi6a8cBCTTTTpaUlnmTAre323YaJSk0K0RF7ayAk5
EItuhySNAYMvsN78T0EDXlw8qXm6g3how1knqDFHSJY3Ywq0obcACd/B0i1zAX2AlZdNBoZk+YdF
kq6dn/7IF05GPQ769+tQ+gEwSlg+jPIkArb/0n5fVllCrL6+WRgiUJvwtIQ7wv/0og0iWFuF6IT+
okzQIwQbywAN/6rEsg3Az4mDCuKQ0z3+S5P84do1kDpnK9UY4jn2kYOCZohhKZ/OE9BRiJLW44PB
omm0NOfhTLDiMjM2v7T21Dp3blcLtGf5/JWkA+rr11lCtRYtz2x+8aoZjJ4r4SILPNgDwcoTw1po
q7ONao3bmcZ/P31KB5y0DHfhTfdDy04lyNdD9u4NKalR0Lsf6EKUJ/dApkPcA5V7jE8y8/l6+Dkf
6DJ519FpPdzj8Ox8w3jUX3hCyIdkIh8IcDkRLqqV65V6w7mZntiqZzn/lz97rAWerV4JvgEf+UOI
wNobyTLfCDo9Qc+1z/zIkPs7D1/AOFLOfs0nqLa4yrIKUAUV8FyJoU5A+2X2A6VNxqlQUNRUGSlx
RxzM4Jz5kthqllZf49BLm9kfjJLRXHOeidSfRH3Xp0ZQ4FMG16NSz2Vx8l3bN6PJPl5UDu0H+153
Lxbi6LPGqWRUhpSqJVlCSz0IS/AIBSTZPmGH3q3mZMm2NCP69hRYJ8hiakuVchoVRMsQGWXttbuK
sdYC/QoCvIwg5hBKx92bB0+z9RMb8zbbL9pvmcEgJIT1J8hiCcm4Jij5O3VWT1G5oxU5GPDhAT51
vBSutvvf9YLP9d05nGeChf53j9JAwSZexVKeXh4pqv0kd77LUiD9cOrKGDdEehKT1Kh5ZN1q/JQM
45E8y2KXwhODZ3NO6XKf+1jus/EDhn76UGXxqbSkjbzCcGyQ4LlbeThtYWDO3GwtwiqWbYbxq4MW
9HJkeCStfZUyL0DVcYqTcPaDohayN2j83PlqcLNMQyd6K1C1bAz4L+Nqd/l29hDhWDhZnrKr2Pis
rgrlv5Hvxsnyfewhh3xq4wq/f1iiu0MOQuu6Ny5qOyVHfce0lbLQa+4yZkMJrmYqVydZtvk9MuXX
ZGy0yeC6rFsBaqCtVMzBadILPjJZCqbxrYLmtDHBhDdv5UHD3yuMtVus/rksI/8SMjH7YRrPUIQD
/CnQBzQmn4TUwAKybUCZ8gXvFAcAZatMuvayrKo2oLPumKzbqjG5kaNufrjlMt5C/NgEPYIhLKQm
rxsSpLSbUhv3kJSpHhP4wqGzplQEUKMhaBop/urlizzkdr0lDYDlijKr1Z0z4TSmHZ9mGTntSZZH
fP5nWoV/oYTnuqUqtOS/pS0eSeL+WfqXQtTZwKYjORNrmJXjj4BUp6UyHu2a1SCeLSfK7OBQ/HZn
h5Y8k+/6M92pL3CVVNVprnvgQtItBdQ1lZseDCIpqdVbshARkuN8NQwsqdOgD50NbwJYzeMbDgsI
SXkSyb6lEQLnyu1l64wy61PVfjd3Tlcgn0meJflSGmtY2sP17G7XF3eFlQ070rTRugIpjvYx0vt9
VGVw/Gu7S8srOe01t+P1/j50NCzgCu3LXkaOVirDO8cr4U8EPUPkh8LohDHHIptZxikDql+qYh6M
9GsRSGRuGtBgfrWjHGvNoaMhiAS4CMGqJn35SKJaMCEXvv9jB5xEAhhAinM3OgNhqQo4IL6HUWo9
CsnGB4zW5/U7WYTn02lK3nQnt8rvyxjPxHqr9XzWSTD+WHVrFaJ3yYvEaQ8ueeJogLbe5Kg8sXIr
DePMPMHg9PvHfJTx/5e/ngTa1ZnNJvEHt6XZwxbQfPggGXNiwOkMHd0tQLgzt820/fpfsfdVEMNw
XG71kHsvi0D+pqT2KMlmSxy0Dbu4J+0smtkNLW0vWyb9szbRgEaWBQGplFzgJiUzPIFOo7y/VHqO
Dy6OgIdsf8uyBq2aLycU62pqBBEDYVSb5ST5DUEalTKyjJZ4kQQCm5IJBPCJr04iOAa66c27P5Ns
eaYt1gDr/rV8ZGgj2yGewko3hNCC0l75SQxx7z4m84DB4kzENPCDNJsqDSln1y+1R1AVUE7k5S8v
jI13c0JRIrtzWlHxbj3RONMf+TZOgSadgrAm8i/8omNWAQlNWYxA0H0aEiQR/AgCo9vlniQnQ9WT
7mOhHM1cMtTfC7nNq2sjB66uWM7kxWlLdg2dx4kAM3AIFjKb5mqPOLK76jFpdQPaH2KqF7Vl3imS
UZVxwFoIZtETzUX5AWzguix7RSnPZ5Qexsyl1OpIPWlcUibcrv6IkGo35kWRodlRyi/KkMEKeJ7J
ea6C9k7zgD18H7B99j3zpHTmR/wUuyDv//DooWIe6aiTzhDPnjmfwJMdMiw9al/mfjH1WZ2zXQH2
aixXAJPcmdVKNcr7NEZt5TN3LDAOQC/OYjIumiS/UBY0eFOS+GztttJRprJx6p9xRwgd45IYCKS5
lDw/zlFdlLlGy/I+ZzYIdmJpRNB90IafU7I2n7z4syEwzlSS+VLHi6idvlAuuYYzq3Z/CgzKtITy
P65X/QAfR2Na/N1+RyBERdArozb3oT6d7ut4nOYTrmz8LodV+8x6CPrM9UkVd9Y96NkRzYDBASSe
Gr2U97T6lTF/+dRCCCMHZktBFie0WmaUgXz6AdppjaMlQpcbVmSaH7OfIEcVMXJlkajU7LDfp7Cc
e4Ld6I+Oazssrs1jVc1VBvVnLTT54ZDWtvRuEkpLwcqGwPZVNJPqcVKp0kDU+Y/7aTJYTvmesi4O
E5r/NFvPCo3NUpYYac0Lg0TSD4Ikr0bZ1A0Pzwz2y1QiJSpZtJ1LQcgODClfrCDv3PmvVM/NxBLy
7byakGfSTzgJ6xnDDsYATHrj30HIGPr+tqt9mG+Yuf8PbSPucyoJa9cnCrBKt1an8Hbqt2VM+tIw
Nt6Xal67LDLa8uKYgOVYJP9PW+3EHizRRV8w7V43aJ9AbbRpwbRumuI+fi5CHL+2PuYdFW5lMTY1
8EqHThN2Xhr4CMfUyQH5WPWGkTcWAz90dpt4YAnBSeI572zdqpz81LeFeFVLdiAzqNs5ut/GGGgu
L6ChaivCBrxpF/jayFPoIeoq5yj8JTC9CZqYcUyr6pJgJF69WTUCAHlRvARaXsmgRykBWGrPIBrb
oBJ5MQvJS5+F7YfIKFrubsrlqURYjGiQEQQXQbM8qtAG86vjterF2BrvEsWskxutJI/irLpjf67H
bWMfHugqyn6NmazkJjmKfG8SDMEIyl7Iu1EujAMLVbVxJCE74+wTBVs3HrPi92p+MwdE984zmU4v
BYY1dGPJ308O43hiDia90LQMswgxu5x7JppsT7x20q6/aNVtZhMYdbIcEucDbHiqYv9N8FPEQAjw
W9e+P59nx28CIu5yZRMfTkVzsdzBPjojzfUEsElRwBWrVRgY6D5UkO0AmyT6kz0prCupK8Ex23qR
XSDW+50EdacIDM19/j/6vFD2STLAwupnioTY8XGg8yNsLYO6QMGOyax88JrmEdkjG4f2QS8EAr/R
7WGBPfT7iNJo6y2gN5NpdBMYhhy5FUr8+BC0j2NRC6P+OuG6LZKRHmHfA6DUyMVxczkPQDUO4bCr
zLILrTeIqmsxumdRARgyn7mPw1Qm8sfMYqoklIHKCmB6DYinFZLjdtOZpwFCQ9TykW2FMOJmClj5
DfzK9pA2uxkhedzwzGGoYOP0W9kTHCEASfGIesgIFZDTHWOlU42Zj98Ibo+qozdCJBGgytWvgc9e
FsAFQWnFjsnVfMnQ+qAh+i0+iHjAhxhDduLOM7b9Ot3b7OfPoXglhu14aw2LgcNoer0M2gczU59c
woTXPxQsSvNe1cqzYApU96CO+yxHNIk8dnsazDYrksQm5Gn7n6pLtOB713Br7UOi8jprClKsCkKm
Yxae0/UR9PhloVyVlI1OJ7AAbTmYLJ0mB6FFQh2C/v+6rRxFyKYwF8+oUTF6jQJ/MqRIjc88OzRz
xsY+vaySgJTR8wcNhHpHzrTWEDrJtMNgxpJdos7weIWau/Z7NV5GUfkvOFkYPtlqRhlBhJvWLOjD
APc5PITQrqhAl1L9S2XEgcXdL9gy8oXcBHw7UnTho9bBQUMXy1yqKf/MvS5sShnbRm4LD5DpyeDn
0IAtRqGvYEq2CYgp+fkeFpa8If56szqkQhcY2SkOSb2P2ZuqFesQksL/Jb2OB5k2iFHFPWhWe04D
yqaE4t+8NDryuXppkkXyf0cy6Nn0X7fvY40UEWZCFrogH0Mwt31ZksNhww0a67W7R3mmmjBWfjPp
2rtdIW7hD9f0KyeS/yOIM3b3FOtvxnfFbwHsgBBNbs9BKW3SlIIWNLLen34oJh8Gs93Xy3uIeZzk
RFBG/xzqEfxEy1cqZJCwKwpgLbXpylRgggZ5X56Bgbxft42hR9s31rOIfHtUDVqV0vn8AP8+1nQq
FWa7X6Eo49AnAOen6WdxAmxLNDlDyX6HC8sNtDoLYfHiIeCI6FNyMMfrQM3kwmtcbv92HHYHtx6P
CstzIZEUZ51zpFZJtFSQAQ7lmCi4rU2v/kukUw2ri+Zcj83m7ynsZ7r1jh/xgIZeSjz1hdl4YPrZ
b3Gh5f3Z0I96NN959oGnVop9wl92KwQDwZBnkf3RfWhjqEuOWb1rFov911I0cffa5NCKOeBJZioL
xhKQ39tlC0GMytzi6LB4UReZmR9JJeyWlfNsB0E6Rnr7d6Ly3X08QkBB37utlLFmV86AX8jyPumR
Z6ThoscwPcVN12YNOgpLFiBoayDgXot+5aUb3Np0vMaSC/XieYVdLQ+YEaH1wOJxuJ46EykCxb5k
OlR8HQoN2yW1XBrYHCoUNeK4nAA41ZS8nJwXsCCsEgffFzZfHAGPa3fQzRIxm7wc7XeA6EH0gse7
kn+T32j/0gwhV4gRusxXXaAwWwf2KtbhH4xgo65DpfjuJh/SKazkt5sKoC2GF8wC+C2D8p+aWppE
IafkqaBm6VwTgSIbKMOYn4kJEUUKconyW56oKD03uCizrGwDZzJXgTycmbbipHEOKlPj+MtCtXwm
f7944rrqrLf7FicHmzzseJEJvoJbRS8KPPZU04Q+DK+WS1pXNf8GZYKFZkhRTTLSYjA2/UMhkuVx
2VERQ2ZRJEFvRZB/JWVP7iw0GesfjxyrsmeoKNEUxrCHaq46d062t8kqfBxkfD69YsvMNGNFvQds
95bHabmhdsosEur4lp1YQKsULx0nSPsvWrqZTSVZKjsQ6z5RH295IdNLi8v1nIXyUR/nCoLP3Smh
bAhUfHDVzNJLloFRfSLCGLo9gBOIZlh8Og9dYh5C4N0x4BY7VQL57Re0Pr/sqqcE6Fh6SNDNim+W
U31uxGkjDX8UXp6I30WpE2h9I4BcFQTnIRY6Vrk4XTCcYBY9F2xRXtrZWcKoyHy68zgxj2Zlcdoh
SRDbC561SOtoVO+eQT1sND3r/DzVCZf+7bhSmdQc+MC3HcHycSbef6Dg6f4NL9xUS0QE0sdQnyBs
WcExkj9J5Q9+QQWdUgzvgPV6tIr6CatNUDxj7JhvoRBpbS1siVYNgGAGgS06fNf1y3VQCd7/kapJ
QaJN9XK++PdIfps0DXtyqjUWJz50TiwMDoQOSqYwDj/14AxKukyKEYepl++5IPqI3kO6wxsq+lC2
D1Yu3q4KXfAiBgau7HcdpHb6xPhQZ48ame+rynsBi3e+Aak0dHdVRPDxtlpxZ0HVY4uKqgDirF1X
78pLsG8kvCqg/B4U6D6G1siETz0vmjZJ88MxouqCxBSXONF0ty8/mKleES/ZVySf6nGES/gJlTak
L1JteLwVMDQI+aSxatl2ZG+Z6XGPOp3yTfaFlIHwVUdXxhimrx5R/VoaNKZiRIa4SiC9L8EbPe3i
4jPOV1I4leFmvi2gS6VLAbB2nJd567fxx9bJxFXwal0TaolTggvpvgKpVUK6f/CphugQFz8sjjvk
Y2GCnnY5/G5hAmfH5o25iVADJ609vScMu7WLPyiJDHY8mne/qyJvXB62GMT/KvMOn8Cdo0NPQNKs
LhPZhKNQu95QBjoIZJZgwfKU9Kidjx5O3P1kkZkDQugfrRBf8VkIr3tlvUaL7JOfAUp1VZrby1ex
vrK5UYa3FyffinufUDbgm5sNvewWFELke3dnXIm4+5LmGmlR514Rinf3T5BEm/6DsVIaRgICqIBd
6i1ys4RYn+bRYq3qF8zj80UGrh/lak276QNUum4JRpo+2cSt4sp1EAoxpJniS0TrrjmNzVCusvHm
15NED/kApSg9YfhMKPc3Fy/n4NAGrA2xQXMiO4ilfxAEjdLOo/8fIzwUYC/h/BhPgZb6LnR57Xaa
+AVFH2RuzQpRWKmzZYB/G2ZjtAgA20G9GCG90NND8xQ2BIAF7vUZqczIXBU4zUxk74FVWEXYuxyH
KdUuxgRNrbTldH2xT4nQiijwmoN2FNMhsqFpzyj8YAW9FImtH/Nqa9hOCmiSTKp5OBe7ZQworg8k
zvxsauXbqFcgFX2AJynOXT2Umwl+cOi7+7gfzolmTjgPPutYZsPq+AdA+KbPRxF5SMhm/XMZnqRB
KOc5CY6NL4wg9Qx2OYREf8ZS2PTWJcYnJY/XF8ChJCvAHNbi6u1jT3BBzN5kz1W0J7pH8MvrvRXI
LDW2JdKwXX3wv4rU+qdl68cN9SFWHMl2q03G4Pu1ous0FvGEBScxewva2m5rFpCDChXSGAkQ1KFk
iUUR7sEAHIPjxfRrj0OCQdCJVSvsQJgMDu2M+Ns0MllAuWp55fJkG+Vr4OE7+gTES3lrsFytXXZI
WZ2/ijiFaZ2DIYT2xW2SHN8JrQKv41sgulyHGdaD2dbevvzXJrZByhGBcJnnt7LC3UBCsBI+yRMb
Inx/t0FFBF38it5CuiEFzhbGQcRh+gDP88nLWIG+yDhgRMmt80uMxzpdPRs7F2MDfSWiZrGjtXWv
sGlfZujG7dR7tQ1SHc6vRQicOgnCY6Hz7MSu5QpY/ZsDrRTJmWQ6Bq7BoZ64hsZvhUJrRUEdNBwK
uHIW4aFuTLDE5daNLiI8JoeHEG8eQ5hdJIA3wmULW2fWSZ03J2zHQcLQrDjmW/NXSAjczYlLSiGG
p9A+/aIpb+gPhmmBajPkdMXBBXIAQ+axiZKjDyLX0VouQRJr8BbUzrb3Y4VDTrFeIJyRSGdByCUw
EMieody1d4EUx/xCnhunw6j0BZMcTb3/9UbpC7eWYKmucypClpbFhUqo3JR7JMFW2+YLZH5BRlob
MFbnVlSg4S2Q/t6k6maq/p439SWNH0r8VxIse51WiJ+P7SgPVP2e5naJtz4mkVYYqRPTRZlOgTcJ
FSsAsMUNz35eTSw9nTEL0+Sh+zJlpd5Ngvz+8IIbixf2sSJVL13kJecW7qQe8YT430DCm0tHwZ56
IZ3va5bQJNrlmfFQFIZTXafXoGC3M4CGApLPWWPPBQ/0dYEWGLflBXVWsXP4LcfJvvE2kBjwlRtQ
74EQLCpMDPcEKYIdea3QF11uYZ6z34vkIyBfrMQFfdcdBhZ3hH0tlnurR3lhBjsOPQXR+hgIInLk
5xlC++rvFblw+Oo2bX3nKU4hJiInQadrJkHJQ22J+45ywIzNY5TWSNGqH1ubUIS0Qc6R3bJflxOX
YcCvQYW6DyJOL+vdbqK+fFWLianywgK8YgE4gSQ/r2NnhfY0zvj+mT6REM+00uf7Hhoh+mb18etf
P9qXrh//LVMpv/i1zcIYQvdKsQQNwiPrvngWucXgVsLbG4kKHDqbVaJPDByCUWEIGwvJqOmI8/u2
bBnyORwbngWATnUzpiy3+U3xFCf/F/F9iZiOsTjOQoqUtCYOBAxT5OH85PdAJRTjMXJ0FJEU4uC7
4xxWD/JOTUBN1PDadEtwaFb5/gaBiQZEDC03YfS0pGVyWb2eXe9X5d0j5jpmdzWaywpqDAcLbv8F
gxjD2eKlqlg7gIxAspzBRj/s9etEUsKLFd+gS4gkSTNx3PLTCTrR7EiVGi7MAIzjrmL+YgoXEcPQ
Y0xF8eZswkpZZBOS/KpHd5FQaj7dJxf+/G5VM/ykznFbk0cvTltlVjpWlnENaSpb74oGg6yslsA3
LL07DeFlRQ1zh1F61IKR2LyJ0/fnDYcdMFm/TRsSRlbkyyFB42u0j3BRukQ/6huA/WIPk1qC486D
xHVRJZ/H/4o1IzLAtflq5KGzbx2cXVCgdSot8+lP3T5MKGY1RZOzCV6+M/zbmOgVEm9AWv8NFe/9
CNSbEro5Ifw4Ep8f6xcWKZzidnnhu9Doj+ioIkd5Egwp6MQWCsaAzTi66R98vHDA/rCS7Kwlhmoj
aCAjz3q4kMN56RbrXbw2o22Tji/7SNZguwVXtmWjBHIXW/F49e800L8doNQHxIiS3fMgJrm4SkBX
8XulzEtyMpEWXYqVdD9AwMWjsidEAwDyvNQu+98r64/yKZNYEFR1zh4mJp7vv5S/XOdx7DS6JObP
qxTXw9nInTwMB5RH6m6OJRPyqU7WBDOpIlVpviVHQBeYoz42P+p2lqj2O3/2PRRyFSMUFxrB6L+W
sxX1dOB+Wxq6sX4a7qR2xoiiXwZs1bVK6oZv3dKmZQfOqmOuKj6hkON0MhvNCt2BfSq+4gQmxtAo
atArhl55dZM+crFdWZ9vt1irHjWxL5b/7BjrzzplGCSrq9R5o3YtxSY13zPU2Q+WRuPFIMhfahVF
jZLF0IzR/sCMGWcvowA8F21t5TKpOX6uf0Im9MpV0Pf0cnCODZP4QvbERwGPIRQfwXemQLzD5g1G
tgdYeHXrgJazipo5Z2piUb/36ztYEhv9c2kIK+CyQB6T/bj1dBZ59wh192BwxHXRrLsyCgVprtdm
nWpbMokDrTuOvO4v5g+Uy6xwnQUX5AuwBiVnECqxTY6b6FPlE9KwZSo2ZRHRtwfF0tGNvGTher1m
h0Ju5Hqo80n6bWclBBH06adVjobFlxDmDOQtenCNUrutSwYn4GJXWYmFS2CGZZekoeeBUuYDhw3a
mFkL+CZSxG2BUlhNPgJeMJyEAz95dZtuqbcwl9JB2BXSpF8u5vTHxndVfQBUHkUOzz7hdMp0let/
aliYX5IXk8oeMOm/MERzDB0vxX2Lfnnlso7J7MUNA5Ib6GduvmmAcaAovxf1g4YG42Ci5Vm3XsUV
OJliP86TyOWerhzUlYrsTLxzv/r48IG1FmAUSh2vYUaEVJIIh/2FnN7Ytw2DBsR6XMhMqcC0TUC9
0ylmUJHieAdqFqbrVwQ2EJMZoqdwuJ2UAJMrkJ+2NdqrDsZbD3//toTlO48f1SGXdYHXqIUfbiGy
/8Sah+PsKdEql/Z3vdTL0kdhUTWqjkmdX9ccX4eKR7CN+xnxZ/mOEaUUFp4rWj3BSwsg3r7ghWNS
YVPAafdK/hPo4jwVTJSNvyf2P5z5girbjKZCAqOpRUeybiJMeK1XVOJ6lxX9RVrUX2cBYkJbd6WR
OVr/IFvXBOIDbiejuM779g2JeZesegKDEN+ACvgbGxRE82XHQsJlAcrLDjGkD+HQk04tkQoOOXA3
kFJ9/Xt9RzbnjRuyo2csfxF/P/j0uf4ONfqZCuDyMBfS1+U759rIbHI622X54TFoO5EjGELzsLmn
kX5eB93hyeC1PozOBttLetvHbcRuPeOD811PSOiRbgipGtavw1GMUzHyy8re6o7b2eI6DtkqyKSB
ai0B27oGAwW7AdDd7yEWcV0dvZ7qVbw1NR5x1dNxrGq4PLqwI2NAKPqCLLBzAgjbW48iF4WdxNYY
gsAeRNptqMgk9WfL4my7WOP2SHpkWz60GCpMHF2/cAIbHfUfnr1Qy5YNYCBXS/KRJZ0cuNkYAX98
84UB4LA4FqMaG2GJ4lj/4IU19+wXB81mnel45AUkQhkEYZabsg2n1jg4FpgLdwqMZf3uCSCiQ0rh
B0MBG4DG4mly/dy3e3g2Lb00FcA78DQy3Bk38ngC0iJ4KaLqmdcemBv2jlVGOYKwCS7vGdlUkTrG
rbosD9kLaMpYFdWoOOINzl+T9EYSSmG1WUUPnnco+tLiljN0mDqvwtw8EAU6Dptguklki3gvo9Vn
oD7ZFAoq6HaRRTeV9D+0muBIvpkZwXgqGKZd8RUd2OMLrHimEP1KTvX4fzaFmDns7U7joGZ2p7N+
GLDi1lz4P9hy6eDzo/9AknF6FJRyZDm//lemv+ukHUE772hDT//+IREx0Tt7wM8kbCd7Dj5czfMy
rRBnyvibvn/mFalINvgd9Jb/yYgSU0L7jaQ7LdVLmyliMmg43rbut8ANFBD3v9zMidgnYPSEnOPL
Zec7o1P3DC0UUz31RBsOUIcZeWTEu/MIFi4zQh33fwz1AHJta5uOdTz+Mag6mMfd8kIqZ5Ks1tYu
2Ipv/bcxuUkA9ssXdfwyF88XaC5CNfVtp+/o/QoLYnoUsIEa37wcAhhaIAcLFv0moKRpMsjzIkMC
4Cuh/flHVKqM9MOQ2mI7xEO8hJOrvuOz1fyYDA9pLlSiWAFXDK9UmV6vyCyQSGtpxaDHXo0lDNpi
uYLEQ7dfpE690jWU1IRyXO44aKF/8FkjrN+GBAUVZ7fNq5GadNPlQKuqIZMsJReHIb65t4hgGdfg
0xGV/ukxkjfk9qKtiWbEQoZfks0+YBYuc4ICZJ1Fa6Bhz6LCWzD1Wtj06NV0YA3SBV0iOv1lJqeh
SKthL+lcBtKdY0LMd91mOv66gwkgkZZcKyUrPJW4QeK093n/hSt+xGnfM4g7nAdCVlAMGut92Odt
DGkjMS+uAP0GhywK7SDB8gOqJEXkQ8c8AHkoSmucjlY7soyh7+ANIeYZBUrhramWZz2OTB6G/bD1
ULjQFlb3bDQv4YIraWL1hcq9i5EMwG+Un4yvb74Lj+++O8H9ix7G5hlV7SQoo5uGWj3zu3bLDwtD
RM6TXjLzoYzym91CftxbLgQZtI+QuYgPK3sk0VWWzV0OZ8P8ntVA0aFEcn8rA2IXNwKklP51AO3y
oi07XKXvNzwU77K/YbCqlnaK6LY0QwjrgWkeJuodTxPPrJygpZxgOuA2V+2L3R3rEW/stq4duTMv
wvB7z0JD8+Skmd2JNhjpAdo+4CGK1W06WhCb556hiVHLCkHoEWWsx3yjIjs32s1fmE1oamdUux9G
CvInTq52a7QAMLU/UV/U80NHOalCUMiThaEyVML6boF+Y6MBeKGGI+3V3rsMG/bI9snkJutt1Wla
buWO9knH9V51bL8ym2SqUfP3NfBbsIBABIjWSesce7qMI6pDewXCXWfZ8ddYReLJM6DLavegdhbx
qmW3LxgFRjHO9e02JTOyF3oSJH0GYu4M9l3w2qF+8LvIdRuVzlrfzOXTVa9+LhJi1DIq8FQlFHE/
oETMz24wNyiwJhqJyHMjDoKp+IUC4xlXi+Tcm4jJc9XC7poVcl3pUnPGUN9RiCgJlerT+0TH3e3Q
uAJ6NphFZHnjIHqWv+uGx7uYlxbqbCJz1RG22RuIiaSNM5vdht9BbcLmbEmz2dfxG7BLhBsQc2rb
WhtVcP0Fi4Fsl+H7bDFwYWPIkod0c/NzirP5QYI+cg0uzHDU8Hxf2y1rtFA00xPzOJtA+QRVQSt3
FyLjQExJ9ETaPIvXqlU3voT5u/HQTr+JpDJwxGbsq/UOme4Tdh9CduCVwYr7BgPQKytMA5I9jYVf
cj+P85dRwaI6Zj8kxImysDdBXl7dNLY+m9L7sqOqC13IP6nsUbpkoduQGLzLZqxq0wIJFBwjsJ/m
Ci3xS+qQyQ3/76hdaawATHMXFoe+t4gaqIYysXt9nCqVBvPGw0OIw9YoI5oUfMxbCmNQOeqgVPNN
/1NzAmVHeHVK12ye5UgiIkochXmrLXctBbKfixRxbHRqIU+0YrokIMh3Y5GK08cbCMlKj9cbJMdi
cfS4JQQdiVlCnGxCSol39TeWHuJZFJ9zVaVY94iZHXXLxuc5sqb4eanPII1P2Alokw==
`protect end_protected
