`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
l8n4wcDTWcEy5LcZ5WY4Mpj4r5ejgBp86hge5z1qBQ1dCLjQxEi/K4P9qBozNBQan1f1CK8Xzgyp
P0lKd0IdIowHVPsK9QXWvOlVh3nza0vSqm3NSQrt99Dnn0sYX9zW5uYDfPo2kuPkbVDHNKN7eIrv
4kMXfwhelRRRP6FX2IvpFQqzDvLdvmdoZr+rkSW07+4pd6Gvmnjza3/HaCGNiZqpncN/Ymue7BKW
scFEeHTP4yOFBLbYgUvucm8ZEAjUnLkj3xEvJBX5KqQ1wmyP5lcprJ7CV1SSbQH2usPeEUTYugAf
UxfAN3b09RKMzBnA25+iaTz5O3f1XKSGjITq+w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Lno+adlmZCO3kbptRY/0Gm3Uf4c/pNXszvVwWAaTZs2qUpEHTUblMGjSmjBwrRnDqU9d+UKYX3T7
09fp2cT123KrncnVGPgDkT0sWudy2AFPEsEuIl1c77sfatp4yHeT8o5H09wZiYvjfcSAGpHDwiwi
Om178YR8fsUBezehIxk=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3i8TgkAkQMB03i7s3ldk1ajR9TtnuX6UNddnIAvyEWRgWgdiWXv5A7S49AfWskPF1ALIhQk+/dvU
aGYzHviYMl1XfXafCxZA6PZMl3IIvWQIhQwCFrpAAa2iMRWX+MjDpe/fVZVW+hqGVhOoTLygn+Xi
oiyp4D3xcmnY/XwCFKg=

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9792)
`protect data_block
M0gR/W8gnex0KStWEd8yS1J1whJvm3RFnjoFGRDtchCiB+wcrkR2J6/yV40lbv/Y6ngOdsRe2TAt
z4qwv8oREfPoBKZk/vtrR8vmzLY2XEVscplzByuTB9GLRX3gI6rJAycBO2SPmL6+7FtzPiYB9xOQ
fSqMOnbnXupyU3BCOkUaGUlzeoaSuD4X2po/QSLilUQFxaOSOJEZwGszHzLK/AeVK8+d3rt7cJol
ecRknpRThC2NOklOeFtDOR8GVIRdr+m4o2Unlu6gFcMx6fgdKGUS+BkBjGbESil/DIUM1xPs3FLt
8aieH+98d+sU2RsxQZKEuBK4UjzfR15gVK6jJj7mzKDTu2gNh8OBk3h6lHW23y86IGNWEs7sgM4e
1YXfvdxQwa0WqLEq75lmT0EbbEMp7AcH3+0EobMqS5KmuASAnsx83LOyqegWA8Yf/Vr3/oGKJ14a
K3Hhu5d/T7r/YOunkuDIIeH7m36S9kGqFWd26rlMTqnGsF0kA9cTGdq8daTz3dAU/BLLiXbGB1VU
0BxmUfzoYXMvVfTXDigSjwOs+a60aEqWbHkeveG/oVV5xegXWApUr9iwyFpuwQetYlPB6RHbZMJt
BMoEdOsgkqs/3AIb4ujYvu7irXxQ4Wj7LkBfw3mhmGevAdTObUGIF0v5l3wNZS/jHsri7TzzBj0r
r5YXfCfRq/mQ873LsxQ8JBU6bR253mhRDCwbGjR/HKbNwIjBrd0G6oTowcRZNWueSe4qy7Drt50G
5qeTkKvUedtUfG7f9FXvPo8px/bWwrahlP/7cQJH8TX6ZeuUFy9v+mCk/Ird65lGpw0/0oa5LShq
0SrfBivpCVRRfOLCNsWwGlsDQzn6vgnB6MMrVe2h0tITGyv5+EqtB9Rwtpam7+1yBpozfdP2SQXS
mrsvRoG5Xi6qqSR8DiqpOWnxZO465l4/Ujpuiu3OjhYTzruRK6De4/TscvHUQ0wOBq3knrdUojSb
/ebn3cwUbonXRqVxZYRn0rMpLKCD3GTk1yfhnWysCntaJpVZS5bFfda0vDXz7N0+2mtTs056TU6a
tAru4X/JGzc1Dejy6sh4rYkw31mFtNbMdpQkOTEvYl54ueGFix+c8/TmdkkL2C/Cj8bybU8vPFG4
g8EKz4xjq/ibZUrvBcxXM5r9HCPU2Z8LmQA9Pn2ZieyF/YiFM7gFOXMEpe/NETu9Kl2WC8edHlX/
6YYkv4AP6o8SWJuXuYZpI6g48tGcjebOc9avx+Hy+020x3O6S2K0xo1WzjcJTxUuAm0+teSLhf0w
VCxTq/8wqZi7QbXHdxylVX9Ayz2zV8Re5naKS0X+7ArI7xYxDIQ4/Yw+aY5xvYBbfWh9ciNWbopf
PdSqCv0LRQ6pnmkWcSS0bEhrr0v70o/xxsDsDDcR4VSL/Fg6gq0ugTibUs44yYH9L+S9Dt7G5Md+
zMpiuzT4Y/hEDiJEa98Ygh6fjuvsOATaJJ8b7evct2ItZUlIfb9xRXC1b2seP9sivNHKF8BiJ0eq
UlgH8bPM1TJGoDFpNbt8jHHpeIX21NKGOipy50754kfh0vKP8A4UXKf45aZwIhIrWgGTCo/KI2cR
03ZqW6sdAAgvShZX/JIWMqdcYHkECg1A9STaKsXsGDh6m3JACdizCNACnpUyaRKjEPjI5E8GQevC
J56XSc3FxoBuWK0TwOn3Su+D86qfAHBcWW9+fRchByBySwY1DjNCO4Fuw71jPOl7+Pu1nPphmiOf
HvZBY/COTy/0mjakWo5uSBCodUPengCuG+phdnvz1UWvQSzCllwROBP6JYNv0tWNbWeCS5nr+q/P
VtSSdZ1iXvzrdNPht6wEcABC5gPTRbRJ5SCgWRgLgUd729CtOdWxXsfsR+iWlUmztjGk8sprAsiZ
knx6qTYQrv2Zx3fx+07ICHSrT5i1/OhSuUER6AE3RrRCVT1/wIvm/1oJL8FRlo1ldV5E9FEZQT1K
XT3wZQ/z1ArcE5bE5a11tKlq/6IltSDZxa1CdKM7Z/GnQMoCgF2LNvB4ELLg5SQtExCR9EZf3waK
KdFuRlJMHzeNoI5marmZIgShcAgcC2sQ48b/5nE6a/QIB15ssENZ/ogH/WYmjoiNuG47tE+52G9T
H1uv+9ps5AKhmdz8lozA+d0QDW1DaoXNSzhri9ADsVO1TmGA8mxR78elWd4ynq2pJCgJVrtPSkEF
yW4TtVHElR53pq5YCDRGg6DrnLNl5qvb9HKDGfiGnnqmOxhfInqxfqiBHO9aAny0Axn46lKi/ZfS
UdVI8STsmjdJsnFDvIHFM3HOD+S5I6oXjzNHRrrbYQBwxEps3H5IzstPY5vVjueOuDDQEfoUb70g
VguIeTFppQKQpw5ZadPFQJmDYgLiBe6bgq1BBLRD/J9E9+2tLSKolKuySgAOHOS1DRVDKbOORZUF
3BHbHKLFZ+4Nk7te/HWAJEIO7kw/A5Melg/6Pe26vEEYex4Alc7WAfgndSad2htwKCB3OJR0VHhf
GZSiBcZEvoLuPhYr6pdxqpaxWKPlGvDZrDr+D0imyV5iWDg0ISFkLc4t+hpGhvH0t6hWsJJJTsKi
s7CJG18BJfir5ocym8V2y61reNLVAU/hHmIa288vnxZbqYKSgAU1Su7bFVkc993ig0r44aUQXrW/
WEbcyGeyrYkpXo1vFjvFTf/SM83xKfJ0SclD4KIUk1HlqwChbQBOFTXiXcM30PfLwfd5NYhzF9wu
7tEgvfUggYh7YbPQXi+ppi2NORmU0//USoeZs/MsalAeD2XDLV2Nf11Sv9K622OlUS/cg5jGuTkg
VvGi3VJs7aT8EAqpf7O6S7CgIyCPl+XPMC3Oj8PagCVpa+bzJTyq3I16G+Yit9O+KBPa+sy+Khvz
Db0SYZCdiapbofH1QMcg13omR5Es5gakylCRdxvuorAZ5q/Z6gh1iwwkqDILOJpnNKTLiRmJ/rhE
hzLEzeVrMV3413NP5hcJ2QoIynLTdoN3Gah/0h+Hg3+JuxLSOGUaTv/VQO24Nk1QMAgULG82x6E4
WCnSGMVvAeoVNHWO/xwZP88ZbzlQvgsGUXNJuiiS2U5yzqlNleOa8IHoH6bMxc1DPPuNhOuozHFH
vPTngS7HDbm8uN7L17/ztIsLlGzSAAPP40KE0RAhY/bpUjE4jKddMgBsrpe2/euXd1N2pycmmT7u
TsbheYMIo1XN3/L/QJXYboPBevLQLjFhMaV4ZwBhcm1pt50ETwWRPzdTNFCoiKM4MNqPcoINLAiA
ub3w9UPVBwIRfWAAlThqbHydv4zATg4UbjEtMwSHA90/FFo19sMZBDgLaUwwO10ywdjgKDE3ePoO
5XlS6QsiGIymQOH46ixz9cSdJXU28wSSUZF9BA0RmRzVPKrvgKAmoE7BAjtYxMLBbEGZAqh+NLaO
+2zfOULG/4E+a8gbbrxRW84OQ1uS5GFz7LFGMLhBWHk1qvVsPePS6JIszEIIGnC1xjjf7y+cuPIL
BIWzu2Z+3uXALEeU5i0K2C+IOHUoENl6OCOmPVr3NO+aYPJnbLsANcS5IjrEeqc0/zsSkRyUkCAC
MdhHVircK5GatK9lpfgzNawm6mDcLzGiak1gTWrQ+KSR3bUILCEHmk0kHCtUcEfZxwwWITZUrNQ5
qTzW/uIvJgTqzZhfhzOy/7stZAHOb++RjlB5kdrJi7f41/KfXhFvZQgA/16BE2K3sueosQjzk18P
2yIjzzBeDpDqAaBrox1GxW8wAM4I0GhbNRsSgUTlXxckZBdugmklbUzbRpEBJBKwvv3r9Kfuu4X6
cfaVAk9UIoyvgQLPj0SAF7UWS2/FIN3jpp8Ydb68dOfV3/I4ij2qLaLLNxNCbc0OxRkRL0uk55T+
dknYx7OeHghrJv80yYaSk5485Ta3V/HRD4zkUfpKhWK+b26uHKp6spSLWCQswPYq+95F/zT16iLw
hDbSyqzCDE9VJszvxTQejOay/hWOFqavVMQWg/5sWr70ECCCAkuKOJ8VCuDIA4DOrgLndhHT6POW
ccAWFB/qEFQ8PP9E5MqVjcf5HcxiYXa5SQUrr7rTINDb1nGzwdYf+u+G2jBvwse3FCH0yIO82+G/
bWDVuyCeFsHhc5gPf1URk92J12senWUuOiUBS7aeJxeAI47l3xm+nvKH0Qpy2ceJ2v3oKn0+SWaz
XBVwy/qDEOoi+0v4LBUgPq2BdqZVDZ1CKBLGZUaL6B9RB177jclw5HCw78cZH2LqU/KNyRoovpzV
ABZk3njPshZqzS0/LwY6OWidj0scHZrmTfVKM4Cy1JVwpCMTb6YoEQrMnr1z7mD0q6xFrwPX6/nD
ZV29vYYAe0LzBkCQZ5Nw02vC9e1pBXHi9/aqybfI9fvkimIZYXnCBBAr/uOIsEyQf/b0IXyjqUca
Ra1KFq2obol+6Ny1+02ZpoOKaGHALH8oU0hj+oBelXM4ruWLKJVaeu/ij4d6Ybuv5f5kMQ5gUPKZ
OHmfNFjKlAg4KBUH4CMjM0uH6o9ELhxpW9RU5z4WiAMc2ezJ8a7gqiHqmyCerS3HNc0kpytlMgBG
mGG/aXR2dKVCFfdoI8fl9OSCI/FjiLhwY55AeEApMIZ9J0SmAPdL950o4DO+4bTphsd0Zmn0KcD1
nRXv6TjpUgFXPNu43IKbL2GTZWV50FoBYB2JLwwyfuRvj4ImEZs1/vhZB6ypDqO1us6BOOPSsmCJ
wCGWMmR58zFWtFmMhhxgEtmaEOJWBvjFwcCStz+8eSWB/jX5lvQZhMSmtaea3tRowAP2raz88c1B
6HhHqEtNp7Z2IMH4PZQ7nlzCcePDCnRVKes0hTqY7g5ba4BS6FvEzJOGOzalWKDbklAY/50ZriAl
A+O9mu02VlSFIluYrXbxDt+yNlERHdCBfvT6tHsBWS2nG9hxmh59LjUAc22NHYk3D0xGFp9m0WPH
fuMm0G/3gfAL0w4fbqfnoJoZDxcuVztFugs4OJOZZpEACPNTdpyxpMQJ2eQr0rjKLbXMpPsZc+xj
VhgziEQtPbUXAiDfAFCBwlHJhTaP+adt0Pz71eW8gt3QNE3PorB/p17T5Y3fmslEiVQWxE27YAv9
fTFaqKQIGaMJupNYSxYiMCPcBCguSBxzydbeddPRubBiOmmB8moahyNoq+YGZ6e6c/1MIdUPZHte
4IYZK1BEBHhBRRYpRI8LmhwxqjlzLAmDbYgC6NK4hfHSYWJGaiNY1Mhk9v1+sKUIu8+2FV0HcjPA
YWs1MAj6WvKPWXYTuMhwZo5hZm+O39eJipbxc3yyIxkwHQvnU8L/Af99+SKjFwCJYYrj3T7BNnJe
mQISgFiU7CkbbMsw/OqGpOW4wekwMG8ha56iSX1Sus3eDul6NGFD8DpmzaSWrbQQQRS+BctFu91X
6jPXXVaFwTYv6hLCz63vutnpQKYeYrX7En0zIuebalAkN9OGzzNZr+BwVMJDKfOPq/MVJusdqk/C
/YEVtADsICsugcYJenuRvLUz09zTfqqGtd3a4oGXi7n9/6c2jDRAhs3Erz9Hivbpl/gIv6M2HGx2
Kkdc1XXMSJ/tDRPbNhobClcRcwr3dpt2yTNAyLaD1kmNjCDIU/Rkwmsx2ptfAC/J0Q008dGuL2dw
//DoWGlLKUBw1Y31Rpv/QWxzumOdt5YoVYiSzBYQVR1A+7SRGQbL8259h+0vsYlyY1kgpfMJCe70
/gSHlxhahbeLRdjjcUB//1xbLwqZRizTJ+zH/XQOfyDAC2vmwsOLnue3ULOKixKELCQrnRTW+3/A
tJziztHKBFMmm/4K4JSc2c9X9ETepPut8ZSqJBHHPFy1DMuKU9zQp+Of9hO8gfmBOLVQIPN9UDY1
L6Sn7coIAXH7iVFLAybwMrCAJqYdChBJwfxTWGRdZhujVcjuoBEuVxaDRxP1j0k9phJFQ9dxBWF9
SEnhjwT0kM8wh6QNYuPSQDFVdi6gao3+duMDFy42yIMgg9FE8O1UppCEZsOQIy1MgSWOLv/rLkSk
Mh0GCXDB5dcyERH80WNFxRjez9a00706JApITnhp3ft8hkReWLRRM1pdsOEbjePZ7ifIWxOXhX1y
X59oNFk3S/f4n3Pah0xNM8w0NUqMrDaKqTigaogxms+2oLjl7SqpIeFD82b2gqhIPba6cfyS7MiG
vKq2RvrL4Lq/xaDtRznvZaOCH6G4iPY8dGkYnNMyRQnpUwbU3f4JK0Daa+hC/tcehddGqpZ4Wfug
vKu5dDId/abGGAwntizpd/difcPoWEpCZp5uQdtCrygqM8F+8PbshBcTKML59/dzjmZLNxDXCpHO
wdhISGcQS47oQrHhqhtxYvLi3ZaR+Yfhi3ULyGo6L5ngEdDrS3PQGa2syfemI0Q7ubQ4HFKDHn6Q
EgBOtqLR49rhUwha9UPAFhAOzlmUx4aJONKnJMVL4FUBiPZ61v//uE3qwwL7VGfKgSGOtpLZ/hXE
mxrKzHZQJIrmsdiAxL0fW+v3VPuocFvTCt4lOBJ4aKms0XOkFCu9yxq1CVnbJAahftLXQvKaycR4
IgIwdXww/YlZnxg6mtkFNmlrvH4gkhvrO5vMow9phX7w2d/6jn5MUwVbolfOAIeYyvqnH3zY639j
KX8ZlOmq3PjJY6DY7xp/N/Ivqqq+J/O58jfMahaO0UQthJi8RNfAsxxKLasuHg9UMZ05ZBfhj64z
cMp4Xf/50AhLk/VTuU7vrDzNtbB+NGTgAg6YD3PCShn8VktLZ6hhtfrOwFSmuxjV7Ce4BpPBrkGu
VUzNYTQtqBmS5h4PWBL+ajBXAzMVuJcRb2zgVIepMB+mlYoQOjQz5CcUQsLkfJc2hMIYIj/Kmqze
aLhGI6A4yeg27B8II02Dvm1ufA5kA+aPBrqCEZLUb0Tj6EaiAths+4w9JIwvR3lkdoZ9adaE6NpE
1wS8TUIJU1FtWFr6QQouGSXVHjqCj81Vcv6nlrZQ7MJYe1iPaVNK2kxLXsP5veZIIt9HgDGimE5K
flfUwlw9ufQyPF1fjXLQZoBkY9KRPHnNmTVrsf/mvQg08RvozKDHQAzaLYGPzyxSeMkA8+2DqNm7
KSIvVgQU2RMaCYK/+rNy3ms9EASTM/zl4Zp/GrhY5YLJnqO/4OpZSyLohsoqjRYRLPWKuUIG+lco
u9huVANqVT59J0wspNGiwcuG/PdNl1d9EPEvA+dhxUlJYhT0GyhMp2HmjjsrhEY3lmW4R3lTXW1m
018FCBpSuvlaegDQJRna5Fbpq5zxsCK1uAhAdyX9bKZ6aXqYubyPVWhCQgPR4OnxQwF7sgnRfqNI
sSxHIW8EDNx3rgI7BdVeR16YOxBnENrMZOBQz9yX92suhsIEDVqRlcNDpUqOska9UKKiOib3uEdg
ZtyZkJmj542q37wnCBhI3ddq7BHVQNrla+uo58sak1hG62+10Z1Ks7YUxcdTGXhNXrda/+vlaAtc
aiUbvGwZzAX4iIjPThCv8ddPb0RlNKqh881vzpTzoM1ggrikGhOp3Wie78CXfeh8eXMgmBwbJugC
+ZOyu2vBOVPP3bRF1qpaGnzBrMlc1xCl6cY2IG2r1gfCL3Iw+DNsWAiy6a/4O3ixKwmK8Rx3OKS2
/3t/grap99efclLXYE5nKYxjMv/572OiczC+1Yh05320UC+ZXW9UfO3zLwVw/vxnyoonRJ/wh7tk
h2WaR6l7zKcW+rWniEOhOQcM/mTPAidui/i8aQR+vgB0AlN+b/AMByt8L+5eLNvMzQeRzpU1tNvL
ubyuxwwI5hgR2FOe831q8qOOwpUvATFC5oew0ujvbail9O0kojMULowekDkjsQbDkYZRVMeiNY6j
kZi8zua4UK4UarySncFFYdQrZuEHI81j2PiyccctMMBFjOh1H5qKqsjTjHpkMKDF+3T7iI5TyJXe
1kzbhHfv+3lwKvUx/+vLu1AvcyeFKK0pMg5qhsPwzWSdwE5bipUw14rro4bn4g7lKuPf8jW/6LFq
zDVVwRNCMbsGBonw6d/peTiByp7qgnNeDBUnUZ5GoJabCsQweSGF8sq22/CMYdw624dAccPgiitg
HiGBPrG4iF9j0kWcmLP1zRbfD4bbYCOa4hY8u/TKDOLwzIp2GW7Kh8nPnwLxLphd+06b/x6gg86d
iEFbJ8enOwom7+rBIj2QB6G3O7G6fJfnlvY+x6wbP6Hlue+C/KA8Hb4IuaSO8pMnMANrf38YTONv
ZZL33ChAtBSZ0LQmPsOYEZCdpdTnlX9AOUWjtMOINku4/cyBLlMFei4kSG7kSqnkFraQ93hPbdMw
iuv+XB/cqSE5rBSYjpWbOIxfgAw7eh29qo5viqoY3HAlqyeu17y4zD9lAcgAyI99aPcudgod27C1
tHV6ZUTPAhPGr/vdgsIbQuY2vsNbki8ePwPXFBBzS7rflgcgp06j2mhmvHqnmQBYC/13Y9OVHnEg
sUngMuO2b6TNmstB347fs9v7O1RhvJsfJkHG0syhYdVA+rgUMV0a6u7/XHqLK5rOdeNvgIhRFdJV
21RA+Cg1Y6LBrKJD+OPYBLHBGHm971DfZlbiUyg0MNHSTuGqz11st3ig8c4mn9jwS5UwXX1GV9bx
Uz31RN6ZANgOk2ZJ9+BVGvnec+0MOUxkmzaoZS4pDhBcjJLyYz+Qoi1xpspP/SMP0HW/CCmnYhRr
ZezDvjwwC4vkcaqIbzptXS/b0xkb3gi6DGa2WAKPpTF/pVIQlTT7pv820hFdaB7NMheMKqXVmMX6
7V+563fBK7QPIQYz8+Q5DdPIkvqB9lmZPgczND8ipPkOF9zQFtZX3GIx3+c6hozfP9QJKSkChdcP
4BrHoFJKjNBis0The8U686Ldh5MJ/e/+6sOBkFZmkgscAFGKH+Oq62k3JEgB8AMdBXtE/vR55Dmu
NJ+XxD6BmvKYJ4LfmXFI1yNGZu/Jzclo8KUEcBxGx5ioT82xMcclfAYjXJ9dorePiRFaTMSz617u
26DDSlF2h1koEg9cKvWxuCRc4Bls9NtVrhivkUOkgFKklufSLRnXj33zgjHzx0gYi7Z+Rf2UnWUo
h9zzMRH+OaJk2tPR5+FydIo+AUXhGiAAcj2l3dDw+sb2jVgL2oUrb2qx5WtbIFVPUBPE5z8MVCVb
JdAnhDDEW64t9yjZR9AbM0ddB+HyvQiK6Z5efRuB9XUTHPCJBKMNxCIy7lNwFKW1eJW/RadmStXw
8DTLUb/1n4F2eMn0U9cXz9StXlFb2/UkolGLZnvVI0e4f1UHpjtK6h902iQLMjsC3B21D3CwPri5
QdSGfHC5Li2R0M1vHsdGMfwl6LvJ4Q/e6chriOIOVanRC8hKny5smerX2v6/LknTOjU8EHITKsOH
o9aLW5VoDV4d2YmmmK4S33illHlm9olv89VsT+q6wnPMOeGXPaS5i/LsI2e3GD56m/UkptXx3mHI
UGlFSXML7Pm8ayQlyPxNaBE3HmcoxAzaAF5QvkwNBm5hcAKUcicxBwrMmvblqli+iHHclQnLEDbV
0g6C1M1mfkGngPlQRYhX/l95oxYXXIGcsFqmaut4ts/DZ/Xyj5uIeV5y8clGatmC1kF4AcUfIVaL
yrTn6XoUPlm7xRivty2feay/y2fdWC6HKjDFErVkylfdBw4O+tFYOWpLdMQ1wPjj8/sPClMDiQHV
nQDIBp6iN3bAopgjGgC88oBlwwe8vH012SPxje1P7bnxM8rP9AW4+p8qmAKRwOn4T26rlJVwA1aQ
MJkEskcxpmguDIrfwcWv0TB7PfDjiPXcxdEDjqzLhsE+HzHgqVhlbzfheZL3u40+j7ItOMepD96I
nG5pRx5Y0ibOIZ81c3ShD4dKq5FRM3ko3Cpar5Y3UYnftase5NqhZitROUrneBQnHwS9BqM+AAyp
vww97Q4qzw02AT+NsAfCdV9KYB3JfKb/AN2Z/T8bzmSUkccqVMBzFG2eMw20oEAD7QAK8wUtkHS7
A3z9FebBy7Xhs+vA+nA82rJlLwRkDPyWVnyjk041l0KVTP/KZUuKAQFNFjwRpVlOAvDXVXCW6x8L
q2PyPmleLPIl+HHMOFeq7Acz2dbqfpjBBmFMoBihYF60ZB/ZuPFE2QbrfVuT5YI6Y4cXCiJeU714
wd89C9sOR9SVxZ5GTMwTuynmQrOwvi2OMZ8nw9hk1nQvHinOzscH/y6MYQndwY45vT/11POMdFrR
ue6jF0ccwrJ6wfPxlnl2E/SYBupXSai8fwxaCyUVEzKBhe/aqHUjinQjHDtSJE7rSw67dwDqG3JQ
KTfwApduDXKDkDxhJ8FSW/h4Tt+XwrwYuVa7rorwlIzkPasze617e5X04NdL4ndTtaAdgIf5YndZ
tcff+w1n0kdeMwXISdNxE3xP/HwURom0riHCQa41S7EnhdwALs0JOjiSVcZwgGVUZgQj1X9XdawJ
M9UjCgAqnJlY6IQHebjk7oHC7fk8xe/VPe9VqNE+aQdq/YH2nIjh6MK/dkA5nF2t7P3MTJFItPig
6NaKGVFQgCJrSfFVQdXBwhvuA6geiWlmbIrcY4zDutKj+v26+WDfPm+Ys5urk5K3mC2uF2VopJUh
hdxdWPLLpluXpzYA2bMHk3u2RLHwHMkR0OGGfkao8DM00jeOAvAGK9Jh8ynWvrkgLkfigCp5we+p
D0mXttdhoaBKhJox9EtMu+5dbKa3bywPDhoz58FeLaiMF5BFH3l+92fXGRon8V6usAkCB9e8Yb0B
RpXA6wghGpw9QajrFM9ubE3BzffCTU+ieaJV/Y35/W2MQus+BjAa7DQZvBE7ij60QDSWU6EyCpz6
DCAbpCRGaLQvDj+CO+RBbsRDZCdpc0sWmxh3JLPkbYbdwbJ1N2zVPM2cfjakB4Gszo6MQTcWZxR9
+q1rZrrIg82vKAys3FFj0B8I4UPZueMXwCtW3JNqwVMkqR9wJkwgVqwvz//+JldhWvAYQ/1/iEAy
w6NbIIy9ELCDI4WJY54EArRjk2nSbOXjK9eluNIJ7jWBcdv7/WixjL2ifFiuL4rCyrJGewqMocWM
J/eh25HiUtak5ilV7GACBhH5D/ZG4ckIIUNvYOSKo2mRf7A4CXnkt1ypvCyiWTK2GTiWMvkVIkql
h7DlBDCSgSkYyHKeBLeEcGwI9dM80ieRvpr88XLgT7m5JJngSFLnNRUedqvxjdeUiyfDYUcdgMQJ
AqPhUKLEH4Z3CyhIUES1UaucFc6WZxn5hbqBTppH9pysuyUm/sHowqpNJmjeMmq2EvULWMlpg7mc
LDx9sC1TutvCLZCf1vw1Kmzz6J6TaiW2sZvPK4WziqUaRfVNQXTXcLB9UjMDU2YjHYH/tIeryp6s
wM/BC0PSzTMTW83zPUQkB68fWQUTv8JwI8wNWTHf50UQGgU2E435lP4q1K35ydHZlM2ErJcU1PT8
yjCeLaAUbkhVDL3ecKN51uEH4UTSQeQ/Vwto1w0DoPRwEy/C1H1MDwTWhq0c3rQSZaH6TV6hKBxd
fbLM5y2kwUGr7UJ8Jc3m35U733YHntGyS3eJG3lwA8R+0oQW8k5Edpb1cw/nseOE1c0bBHYHjcKq
PllQ7tJXxsKbmnRvvL9y10jr7zQYo3n32+GqWLa7J+EUQZGsuTCuonMteNbfJuAQzWZTX45ydSjj
J9IB9GkssB7xBtfd8TnD911+mu9uTpjbXIGoTUnUGlfjSYJa/qeGJAV6WS/ebxyB23eYLem9szfJ
LmBOSfih14M7QlQE/sY2DWd/YEAw5+wMTg0cE7XxjKaCKTwBFxWghjCTCYra99bt53GHghT3ust1
FVqV2S/yh2Ho2gVRYEzRyecNTA10Kwt+vNW2Mgspha58QahLxlbFLOJUNnKA+XMDjAeEzrDAVlYq
FRXqvJS/HpmUxzz1/I791GWwSu+JMNZGHMRF4B6WfVCjKPL8X52otpO++qXwTbWLYgIirHA0QwEL
KaDsQHLzmpjK1BT8j9kiUqjJGvEAbUYfXcInd6L3mLOE0RPJHy1FiQR1UB7QZTJt8JmtUuD01DI4
BP677huayCHWJof34AAfosIGooaquEIwFbC0VWJbLzZzyPVwS2B+D0cvsCk9Gu65l8nFa0FPPoOg
U6bsvbhL6TXHfCPN4ZavJNPGVrloKNCThZ9QbgjnSgKQNAwZpPjusaosQ/29dPVtzswpdsrOvczS
B086B1dXEwBWxh8T4jnvBHw0R6GPrkcP7nWenznmhCM09MPTLgYkMWJ+RET3/kY+onsi0MI2cB25
tHnGnrDzb7QZ2fkKImD6v6Oe2m03FQcc/zLi7CywCPmmKtuyuWWB8TGuzGn/5lmfApOfz9ENJeFA
99Lqv1GiTMVRuRZQTGwsscphylOS87FFKK6PA/I81WHwSAtKr+7+DM7IrjrWQqtcuitDdO4eBdbN
QITwR0rRvT7CxCam5Himv74woWYStbx35Jw0kY60cyOgij0S6l/cSBEJcKBhEMMZdX1/XBgjkg7X
lxu/EqPTFyp7zpK6BVpfth9LovLsX1/KngtZGKaKDsU17q8zX9hgOOdiFm+6re3cVPRYlPYEdUJI
Lk2uibx96u43/ubkMYIDViLr4TCLbHTk7vYSSdGVaU4SF1xVJ5sqaxiIU1DPzddmicrfuRqLh1Au
WvYelm9791LUWkUqsNnUUBVK5uSub/m/z662+BPC/SNIe2qo3hi4pnNawPYt/1jGw2zyIf/Clo0p
KL/fKzXI7qfNEuMMhaN8sWV4sOQG9x9TxiXxgV/PRRhHEJumssSxWOotnGv8C4VEoeW21KYlr2WC
Q0rRsR5NrhmeygASP2c9VwPp7u4T7abpFODfh2kgtPL4v9FBYSsrV8j6vYeY8sLznnfejwxa/S5a
KHENwRr1bPpQdI5gMn0gBs08gKg60CR2OkzgZLe4efyT5rh7LNo0zIQGlQnT4ZGn91Oub46ez8LN
pJIZxCApaDT4lvthsIoRCmcgbq/CMXrNmeqTS53njiWzeQwpraaNyodO7NbRLfJW4vrpMfiQUIN+
EuEMw697alzmdTk6Fysic7YmYKMcT2PuznPRQ83QoWB3dZdpXikB6yAGk2JX
`protect end_protected
