`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
H8ZfzHjdLzSHJmRBkjrFH3fZqlwreqzatCmAZvV9VgF25Uqv0AhftISV1PqhWmngK5DoZsNcGs1b
7Qw4nvBzHpj50PHJiooaw83IVz9guLK1njTFkbjvngOs3FgruoIUUCnlgxknygw38lD4r70tW/bg
9cbP+y0I3PFwhmpAvybndDlqNC2Si2JRsvGPVitKQoy1eFfSmQA+6u6IYC78595SYX+qiQQG1p4b
qzgkMpA6+LlXXr0nzVvam/ZGgLyssmWTruDpCQvmVF8Cb7Hr77y/hH/MC6JNHeJLmIv8BjQo/+Cd
DEzLBYMU0DEF4k6Gg1kW7wEVvQ+CaglpkrjExw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XhfIs4HN95yJzY4E0vhZvmDfsGFPVOGU26SJjsEHr3IJEijCDqWxUowj38d6PiVxsv8khh9/pU+I
wIlXe1jVh7FOMV+/bDJxiDEwKWmNmD6nEY6POGgY5G+5etSulvVAK7aap1YCR3dapiN05TE0/sQV
YFy8frUr8b8yaWhMYwI=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
s9tTf9LD0xzM4/iWVL4fFSdgLO7HeKVOuc1BXfvXj+fj/l5KBvKTQMrslz8Ko9PKNzBoCw2mLgl3
0VluLneRQW2ctwd/ABshLyDCt37qbCHqjQRXHnqAWIvF7ehZziXsLo494LuU4QsadyIqtOZl8znr
bG3UPmI4Dk66UaJqlSE=

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16816)
`protect data_block
/u3yPtsg94iTgK9JeatCHGW1+CLn9xjNkmE43p67sX9aGkpAwRX+BBBZtD6z/Q2+U78EMb15Dk0f
d/JGGmqgXFUO4vynpZgGcwY9gdN5KdbjupdwZofHww7mo43IR7E1WeyrJymcL/kv7chlQDLMcVPo
3e3kb7W0Evom04hqG0KWODPdZ9OjyOOe0VT4TLT7Vf0WYOxr1gduDDXCU0KPt0idbMLAYNR1SV92
ZS/GmZv4rCbuxX6swd5SYNowTuwWLcqovdYuTFAjeANVPflEroRDxDi3Oli5JzjSHS2DyqcWPWDC
Cuoy1nbL7CTrkHwBOzRkmABi+VU8sIqWvjFD+U0VbiN2XF8t8ZZmIeivpABMNPZHnx6MU8eaCMxM
0K4W6eIUDLtdi4LXARiQUrED3wmYPpJZIW99IFWbTL0tsCCaOsbV1SBfkGQGyl4cY6ZqNbP9qUHQ
u9H4PCzoE3EmckT0w/U/uST/6h9wl3Cl40Qh9K5ECknNX8aFXKJI9hS9qqO2XZh1hTRJZ/W3MN7n
vlXe34o1CbUWI1RIhI+6F8LtKEMyo99Cze/LaZ0bb+BFEXUS3l/IYf7bDWNhJw5zKHCwLJSIqZeD
aXaIxhumx/mM89aWYDUNgn/0eTmrk+vcxOA3wF1lhMdle0iuKEtoOkd+RdHHboPTANw3OA1qSWO+
dIhB8H6+0PL2FplFTsNyWtWFKfolpFMzMlkXX62w3CJaKyZkSvSgQhs3krZbYq99uOENq0N15FyL
q4ybR1B4UhAsVp3MqpITgENsitVIp/EUJa//+IhRiv9UzOzSluIzxBI4dPfaHqB6TzAaMmKUhU6V
2Lo7+4dxBWKaWTV0E6+3LWtUVnkXWrpDv6rPxiTF9Va+9gtq1EQ9pRQcKsuky8VqaeFGONi7P4Ek
FzeAo0Sjo2kKff8n1BCN8fLso40DZxLdzVWRr3w9YbJpu/TorpU3GsDb6fqm07VT+ODirLEtv4Ew
WQK+YwIbrQmgCtGO6X5gVv/XKx7FA2lrajDFw/SG3ikE1NPKyM1X3u8dLmbzucTo9RLilBr+iPsy
Pn8qPF+raNJncEmrIgFHfSyTy6F/cO0hMxhIR0XzMMtsM1aIgwZh1LWgsr3Y81XZqKAQzt6RgCxF
a1AZjMIH2iWt/AfREyn6uwOU0MYIyl8PF0ugLSOL8U1S3+Y91is8pAkipF5oEWhbKlt8gIOp7gkJ
aO+c5MLZwwBnNOD1Dpzmr9fjzetOgpjpQWu1Puuxcw4395cTHF+jTf2lYOIRA3EvVrFx+HGfHrYU
37njBfJU/tojiH9CGMfwjtv3XYn+dv/1Ja+Ky5L36BgxizeWugHimoEP0mo276EgTrsgI/RIIU2M
w8+SLcYyzAIHTYiVjFFovJ37lHCwP/O9WMPPUYNQ4/hrG0cQzgMIGKzo3EGBr33SxPlImCbk1z5+
0cgsSDhLYuCeyTu0N/mKxYYI2+gp5O68GDhqY4YwHeT2ThQ/LXzCtKwLHBQfx2K+W8aeSfkSJRSU
+0b6hW5UtbFTxpOUYFZ5Y22aMijGff76Hc5yMI8DHCMoPT37mUkzgbLL9Vf7h7x5YRAnkZwFZr+O
m3fBfja/tEApPgZ0+FrizpVZEh13893/OtFwazIYP9ePWExCCHiZ3EEUQVD1PVwOdLkMh4rBnAas
AiMcSwRq/Z58W12m8mzpeDQpYT4z/fLtE1vzJkJS1GyrzsOAzI30yU5BXkj7RwmLS9I+1n7hG3Nu
bWJZqvNcg1eGZbkXrgBizFURp/49wOnekG+S6XF0/mXT8ESRjHOkccxJul/dTBOXh/qB0r0hUcOH
GD+mJZfHrPE6YTetKYxI98mn6TLnEnEMK1yW+980sq673W2JaZGYIB2vimIY/UtuLwfuIOEvg9kV
A2P4R/mf2fQkmL0AvLD8xwHdcZ7poFaoGpExIiafjsy/t1LzJdwzxOEsM55gK3poeAHWB8dPmCQD
4nTZ2bdo4UNO26+8lFAY2bZbSs6Fw8ib1r6a7MsVmbHAqcgItdDF3xQf9xIjqYz+xALcv9g1+N6n
qsrWjcfqu1wUXA3hEXv/ySXUUIByoiF1fuHjZpI0TLR5nXXlcY0h2L0Xb0flPTkt2Pc9dc5eiKFV
rU9LXUCIQTgXJQlgZJIfFtm7YxkSUC8dLdTSb9UYSVYqWs5WowVjA81o8ltx6F2mPOSQvUiZLRDs
Zbp32wFTYDg28VyWPxzg3IujLQGhmcm+4/QkNb1/oCUHd5vta7Cb0QT4AYXVi5ueXESA3BsNlQOv
1IqvIZ7obNJ6r4KA2RVSKlE+/sA6maUar0aR5mArWF9nPtw4deePEScne5vmrcsGB31wk7hxeG3C
SnPMUN28vG0Y6djCf/N3kS1Z2WyMC3GDh3/gDkW378DJ3o0KbSm0bM/LuCol68scFqSR7ccxISGR
pvTi/4xqetIok/pWAQDubzRy7Gs0YcxGYCANHD3tDwtIzpzCKYJ3VVxY0XC/3z8Eny6ER3udMnZL
5eVAyP9evPgJmuRCh3eDogquOHMmyOoUf5hxS39sgXjsJ5jAW0hbRzZGiB6PGWReYj59BPv6UkVW
8PxLs7BpiBTFUDRQa7V6RdDtJ6rVjJe6U0NjGxl+20QVtBTBNLFl3jaFy+64ri7sDW4qUAQzcY5j
Qw275+yWuIZpBDd1DoSTW4LQvmzzG2ufwyWXXJuw61LWFO8iwBtoGz/6XdAcrkyZclNtyGw7KF3H
gAioe1NSnpyASDy0ykY7dBt2MSji1aBO6qd8noCdpSnkmMsuJCn3e40m9yJPcuGOW+kXCOkTp8xf
T2vAq8NzQqiO43HIPk3youCM8BAsQteUWXCdP5VohDhz1exHd+YxThW77+jWesdRAAxq9xkxY2Qc
TXSPLkhKRCPvIEN0fJ2v1Mje1NufNf9U1NJrU6zi0cipOlKUrVfsKw8OOjU8SUKdJfO50JwjMkxU
kVFQaLAjdC+2vVWRBD36lyBUVjySodMeAppk2wdciuc0IsMPPqXLbnVu/8qxfGL89lhgtEJ6IfF3
xSVUbajKcuvhUg3rLUh98MGhkV7ELPskUCoNr+eTpZ+91p9ZtwrG11xUJeJ2geKv+VGnSvtWQuiU
ti8n/csltLBkORGcfFqtlNIxiAU9Pk5y3nB7rsmgBI+D3sgR9515SxkuuuXeRwv6CIlkE+schs1U
/9+O73iE+9KcLBEjenYZifn03gVlKCa7CS7Wt64OVe/I1KWSHBhU9hQmvSKFZiISY9dY2A7Z7gZQ
XRlRt046HgdqqasW4warWFBucums4IAuhWlA+MXtAqdgb+0jyigQBXTyJNxAv7+D1EI5fXZ/FBS6
lpu6DSM6UkmsCQym+ho3dOhrW6SjIhVttXeJIFby31D11cVVrEj326N2PTOY7N0s3plT7kusBfwK
RTJt5lFJVkGI/BS9c4K0CKkedj79vf/C5qlbQKEpscntLNtq0ex7zboXaIbDfp+NGNP3YJLNXaP1
HVP2VlBjFQyMWWblqFK1ESggB18xNdtNDE1up5nSoODDeLN27rMB8amfYOmoKYfq2dmU47zl6FyD
NdynFn+nwecmlZzVugrqgMU2epdcmL+capqhT7B24S9t+q5fpHH0VMzYkMSpjS5gVktRXGxq+ZG7
M75oY/ErQi3lIVr9qM4vt95Q+6SmUgHXBYlFTsFkv4m6qtzPCgquGjopdn5bfc3zjzr60ymCvu5l
6R2JbAJNyyaxLRQ9LqWGQKp+eOWLHLo1mSEG08EvQy9eg5PmH2fyVqfwLmsdWIgBFwbK/kjHmazj
V0aDdgj3qMgA0BD6NZw4i3gVfJ0bRVzEe2QDSYIQSux/IcAujEAo7nzaG/cZ4PVw8KiihkfSQerZ
bHX7VFpK5lNpdF9dH8cA4BDZwQQ+QT0QhbsVk6hrRJbHDhJGzMVefN1L7+mXPSH3G66L7Dchf0d9
yRXtSCCwQP76qtVYwWEm9uSI08L+bl4roW72LHZK+3PeWoNQXcancAb7DLjQCfmFwJimmPXjc/M5
Ms8vtrnpdEpLv1B/SLZi3m0taJauUX/JW60xg0vHiijXhQXfgnIobHHrmuGttKWSnOJm2f7vAyhR
RSlWmYisNqd4wrRv+0ZUeRldgZhmH2nwqge7jRtAbPLSpOdED6M+odj20+5VsU3nuDvI0DlYiK6S
hgYX8rmi1V7fFSHw44CqS98C3GI/WKCxjggBGGuOrnvECM0uzRQ3Iyk5YR2cTA8fH0OOF+jlOyYD
CXobo4kxz0KlS0CDhotScsPC+X+bM1JZdCjRM4oBTdS89Pw/Wqx3mGgoLYik+Q//450QjXkCzOQz
RrFFSU682WMTAZu2E6BdZmTU7gyXFSD4Gc7PZRVPI1/SEgJBXMgpmHXLzKwiimqt1wVpeYTW8hdG
WAgj+VqHf/AnvLwDS35fQnGiXw5rZBLcl7FZ8LAFrf9Fr3IundlSF+IJ2Sbx0DhL++ve1FMJksVI
6PJAWlQkY/CME0Ot2DWxWpjq5d2v0nKjOpBDyhihK2c6fWsdjbOMc94qTVrCOTlfzGlyJ/ccW8ft
XI50BcyohQnsZIDrOjUfqs1BlctcnKdZYvEFU9rUFzSf2frz+ivsJ7SoPOpuqtG7YnkcAb1fW7ap
2HN1ThOUzhVbNSazkvwNzAUUbxmR1VzsOe5djWmZsxqWf1iMgPHjoin03FHkI6sTOVzdb7MSyLjP
VhH5vFb13vSJp7wkdnUlC6Hpgo/7xgytO+FhqrKeWj6QYCFk2qssbVKyml8HkBm5nXPnIpbzo8pF
FLAX5d5MFLiNiqENys8hBThvObxa+rvsfAihJmvHLaqAeMVJa0YAImhzbGsFtWTgDRlScqdEUrkN
nnOZWTH5YNQjN5Eb+DNSNk8OGlKCxyxxXF2wPTbSUIEZL+bsSkgjAL2/J/mxPzyAlTNYZvofY6UR
Y348bGqtBSleTD3ykM8L2b9SfNXOXJel63Jmo5UvS/uWyDbGPrFmwK5eKXyc40NQkrzrhAEmZlCr
tRZETpywQEOVr0FjMVJOwT8bKzwVqL1yEVt7zVuIE7C/A8u4HFoOucVVRUBOVhCbeCwUhA1aqeAo
a2ZHeVrR2na6nZ8sNdxddGtLrTgJsp/He8X9MXdSq/DJKhPKaZ0sWyVgEeLfHjxtYrKERGzSC179
PVFqnOfSmwGNZueoie3vd+hkSYtE72shHsIVvxHL869RYPbeHHLd4NS8Z0JlcvsS9ouVWudkjCor
tbvlT/+8c7X+g/X76CUF45qH84LMzL258ZFJFBFBydqQL4d93ZS2CR+Z9A9jULpgXSlbCFeKNVS5
Zxt5XCKVJqAfNOOyYnRUOb4BBnnsSTq9tgmgm+mrilkzDDVc4H38//eFQ16IkOdXTb9F0NDWR3T8
tRD3RLzUYWKv1LqztwTcwsrmQB7cgpwfvqWKBSGvEJAx2Q1WbxwUSRKyri1WuaRan0g65Kb7tnbU
1w0ByXfBG+n8R4Dq/X21Cz8H45qVNa/Mqjx5C6Ow7O0UwvTlLmdYZ0pQoxM4erdSCx8i1gsn9VfF
Gmiu9djX2cAbObUesE7xxKglu3SMCrakGIEIz5UDA8ElrZCKvD1IiC7iRe6OnuaqYVenYT+1WLwM
L3bUg6+nk8Yx1BkecQKdLwXtlgFeJH1PuVOmghZFhYGc/BYFMJ01JlvjDfTIXsgFSYL9KLNzXHdY
+dx0bpbC2sX7vePx8DUo6e4+A6PqvT8EipBcVt/rTJf4fa5CnFo6ThH0HVpXpx2HdKNrBjA2aPM6
Wn29UXclbRKDnsvO2cz0vAUAsaJkpudSoy6HwOyP3bG5so9MzpSDBjrKWb5x+TrsMcdYTsLUFsKq
xNSt2h+eSWr4O8IcKNHAnQ+np1UgVufhVk4mViamNDSKLNsD0BDPmGE7E2+pKIVN90s+o4XTf+lv
WWZvtoBqG6wmV1FMsATj3MOfQNyRYW3qajmGsKGD/8fY1gAr0PhciOnLa1/eA6INx6t0uLSZXGa9
Yu0YbTj2RwxRkMG2JyRizJrgdNwq713Ps/5iTaXuyQwpmOhsud2bcbvLVnGtCM4esRlY4xym0bLq
aW1ANzkzLP+1+XVUzOuph1jjXB9HuhM+CMgXrREWgAjTamZlYRVJxBcb+J6Pzta7UHayswHjAaLl
TFFS61U3b/Rl3cmNxw/uezLkWtelWD0X3jSsNTdK9GpKAuvOkEnPIsaSkgx8xHxJRa4Z577ERXBM
Sp3Uxt+MHQtz0YJ3L20y/uKq2ojuCs7esV23v7sGNFThDke+WSxdCBOKB8HPvzEhbyAUOEwT4WT2
t9E1mOO4nVKmqDvBp79g5IA3DenXlwIHp5k0QnlAGzbFaIr2pkoEh7CoWv8l6SKUG+bEqwfIkEaV
OCmpIlSUJk/S55vhzx+qKcIyCG71tNOi7URs/mf89AhPY9wEgedoCEWspW+WVqEZf44cE8uYe88V
6zS65xHICrKPENtu3xaM08iAWFuiblqn6SfBs145PCwumEUsi713bo0MhprDp12/pjS+KItAwmQ5
nHH2EMTWhFpdmTMut6H39orkpj18fC5mzmUY+woAi144o2qJvGcuxBJKGnkzAe1ZlzkV96PkPpzL
kQKsZjWXfWL3D2392Pyx+bkR1ZYVhii6yZkKCPdJJN0nwIMkwoPXdKBlr2nrQKjAYTFQaXiD32Rh
jv7XlJyXxKz1whPXkCQCQjckJzX0PbWrZEOrUG20eOXwh9J2ZC3AdjYy8pQdVxmXvWVdj8CwinCI
P3IgWaZNj+XU1mrFcYKGi/kw4J/kVb/syPBRSTyiPssbyIWTTzxoQev3VwLnYEsDYSqDPzB3wyrK
bb1huJBR/+7bGaMOuoBxX7WY3F45hhrlvWgdEA3iTY4mi+Zec4YXSFqcNuMP/q0I7t/rbrrpC3Yr
wM3Bs27ZTR5Iac6k0AGiHqLPN9XuU1qZwig2gf2OAou6WWEGfgX1DpvpqnXh02NOEbHpS7HsPKV9
uTdD9anXbqzbiadjjf+EJmhtb4I9gH4GiKcIhqEfB0vjtRUJfEGh7v+BVPHRXnkttFwj9QgwuG71
pEbo/doRFiIS9WM8U/Al4kCFUFBrIlpHD8WeP88C14qfJefRjpjnu1tJ8kswdIeTeJwqHDudfTmd
5mhb9dMIopvceAtI0VhM7q/cn+KF50id1I4mRXeVh1fVzuRszBunnuzsVF2lGY823XTA5a6spunk
ra9PjgMsc9WO32R7MQP1bjKyJtLdygSvP/LlbyfVU+ZzoRmNX3HBSBnfFi/xsocIa9YBrIJGBzuj
fa8+D2G+YzujkVvpW5nwRCMQGajCZmbyiox2Ozh/a2S9+1KB4N0ft6xFYi0umCzhZ800GWz0nlA2
dei0jGJPvlxrjzusrjfgvNQlxDpe8nSsCHb0YtPifZxjezq4xtmxPTrH6KoSoBddC1zDv4MD8umc
BqMQcDOKIMI/iT/zp+kmmjUjmzxo9M7hRG0rBnElmPhONXGdkryYIYYkl0Ioh5LDtEZ9oPJCi0f7
najscX4r7div3VUHXdI436rFcqhpj5VuQ19v1Low1KhPDL4Y4+aP1xJpgNpzwMl3C3lAa36UFn/c
lA5VygaldZ6+FEZJydwm7tBGccYkZi5D3NaAYyEeUTAk6auj1kwnOyrA4bjlKzHJ7HaO22IeTefM
fdfEImdXr3MTyw6fI4kGYY/CCsiEaY29U3NwNrWb4E1EoftcEwAgpHIbzYl3CnffsOROTifqnIvi
9fPlnURbfeByXPAz21FaPy4q0zYHcs9Wwu+vJgoPDSTAB2pN3GWGMh8fYlKBv8Rnm9XYO3XRnrdr
cHoNZHy9UHEmo7JDaizWGIRrreWgqEu4N8utzHy/4MMo4ZtpZk8Iwl/E5OJRKrZXyPgCpscmAJrX
+3oY9l9fNbT8q98goNnHiGmobpawRNfGKlY+X3VnnVsZ2uaLKvcDdcO6AHnTlyLXSpG8O2dzp3cA
mz9xE4YFUSSOxF64mnWHhKoibE8YvDgp1GdsYXAR8cgj5urtGxuQUNouUYzSWA2GczNX7CdNcV1G
ESmv0U+fOne/AQShUeme5t0PqW6y+tW2gtxM4ge9kUJZjWN/T9f4HC3FEZgSLqF8MG31MXG3SuEX
4j1i4ydbgqEgjXRNlqiQup+izu0p7r5WSJSUWUgSrbdIvD6s6tAFtF+BLoL+RZ55wu198/HA0pzX
8pcP66SQzsReg+vOnI1FBqewyyWoLfjA8HROafZq96NzoYWhUPApdBG8d62YYVS6aEbvEai8O3OI
V1vf/Tw5pwdo5yAmpS55/XOvub3uObGhSxTEHLdEIcyv64FAcLy5Rxg8aenOBtYEtH+j6/5MwEsA
a64123q53noDeanJ3R7PjIgXtrWqk3caRR5cM7Bv7G2C1rHt9u33+zogSYc/TwDE4B+xtmG7NfNJ
xyMsh5R5v0WY2lT8CYsCOGKuEkrQhznFRjZmgUcrC/WUJvZZyD1I7A5D2L/UI3mLx9wHV2bwjXSM
KxHxQtdiPR9m65prlkw8+G9eiWpwhwz/nhOtcwRASQajaUptmKp3dgGi7INFA+MBfnCRLM4Uq6Xw
2HTi4eikJ9YD8TwCQyYxHd2AqMqPnsSYk0ihWLwgHFpNuvWEA9GcnUeHe70zfav7BMOsnMbi3RJd
1qDAQyL2ZoRWcgToxpuWpGT/zSFKK/5FPP8UO1SX+MlpTdbqx4NN27o4Sbj9Bl0mficflhFhiS9F
36UxHIcfFEY9R+NCU5AARCQsysUe87IVI3UvMckXLG/zoRU5YMRhyDQJtP03F25PqSrd9pLmxD/z
koGpuPM6GMv84ANpPNpux7IbshTnE65Pukovo/uZv0fr774azMcUW/INnOit2h8Enuc3OmsigcUy
1HbPp7nPFyB6WioSDwbG53GgDwVNwAlwYUE1WnLcyZ7U2LBmrZ9OpVCiJkS8nvLyAZ8vCIyUZsVF
NsquJq90WAz/1MlPs5vDkQQ4DsyAGJNjSZ6NZLExoRZWVcv4FJ3qBsGmidnL6CXo01U/jD2OTdCJ
3Rb2K6S9od9vIaiSkBiZ3WaWNgkgqLSG7f2ueXpNxuzHevlS0N9HC7Ml8DoMkiiUgT+jkY2Kzx5l
amV5gEEkXB8TXvA0Ad7i2CChBAbHo5zGNklf/Biuhz2KEdt6LnxY0KlSBQwhXeeL0+MeRPPDHa3Z
i1Zk9cYRJ6sNqmU5IfjQTTgqkABlxmLUiphmkvji32wkFYXRD0mZud4DHPGf7DO0QxVla5Ctcec5
cq3+Ns/6zyrCecD8Qdi+JKoeIIITn+NeoTRIRiURgtjQVI8QwUNzdfTKau6fAlnFs+AFCQd5EeFl
s0Uw4E0EEsDfSEUfhw77npx/Tmg9d7A2wytNBpRNuc28Wc1gwBcQom16EWB6qgcSdTMM44Lpkucf
VmrrjNCLsGYMk8AFcJS5WCHMUNOiubrX/leGbReKj96KOg04IeBUXyDI8NL+UQppQPvYBu9cjPPK
72FfdyXHcHfTNUHmiprcfDVUXFmLKbM9HekixgVQGX8slxTbYsQx1roTKD7ix0UIhCE1PFRAqgHG
r9dNwPqrhgqTE4WvAKRMjt7LzvGsEQv9dGwZU14LMHyjWfP0q+b7xin5hNeX+JRH+y2pNRtPfIJj
MSK96W9pHISS8dmeVMHN1nwBiIym3HZFBkzv58hzZWU9+SkER60WJYqghPlXvkvj2/h7G4Sdm4/r
2qlq0gj2tI2w8G2p7mX2oc9nWKMvoFaM3kAqza0iNRN51VY/u/Z9MMUJ7qmUo0NEO9o+4svLCi2p
0G+ziTUsh9bVmZjWOeCmAG9w4Fp52QRN69PbZGipfRXbO3ohkmMfi6i0zzTW7kj0TjnavT+JmPSq
Dp/8jvyyVqcw9aqlj6Ale5PtPnmg5tqYAnE7ll2NbGzzZi7MF5KdSYnOfbkg2DSnwPIRHDX9Ir+a
tNCeQJsQHmY7xlGhzAPDRqaEn/y1W9pNoKDCTgCpTnaVEj5q5h2s7FjmZgXHZ3KauXaJQG2YGjKM
/HEbrZYmp0DZ4IpWl+fUY5nwndgmfU2g1ABIdXHMc2EJ11HvXGWVkOfhy1kjx2OEav5xXSGVJ4oX
VKCycn9kI5BNlEQS1rr2YcLeQjRBosRfdN9k+QaQbHeVjPTQ4lhLLoFd5dnzM6AiCMOp6YsreKh0
H44IAx71aOfhIZGUkcTFe0sxVckSxprFnN6dKEACAj0DcfyydlBvu4ICjEDW0vto6RsQ71hVDYOf
lj8cMSdV9jL1a674E9X7ZQWZRyIT7i/P9eIbGuD1kKm3WfE8uFVUTsBhQ8J5PvNKc7xxsBQu04Gi
WbZfZVtSU99Optcm4z1PudeTkBzZ0SbRwK9bO+bcTAdlo4TrUz39zu+EnpjgV5DBwka1brYgg/4u
CpW0EZ3fTPEz50/f2VO5K+J1U45uMwjZc+TyKS5n8rk96L0fBaSztKflJqGuetdaTBZynbGGiwFW
/q5T2GfADWM+Yp0CwQ0E4oQ4kor6fLy9n+6PuwfcCZa0j8mojVt/0tUCQhFoYCVllqC+t09bWw5S
1GdViWYRbz6VG1CI4Ovo1l3gMQFu4tuPZ140XJRqiGmzaWKvScIq3AF17QTtBCHApN3tCswSiz64
FUTtmapGlFhk0vQ38vWHvkPZQmGWz0VrdQcLy6s6MEPi1gev8HKxRyi1d+cbvYC3Xd3d77w1cGPb
VnsmAWuqNGMDfkbNYsAOwWxiV0oICiTJQjD7eRVkZO51+B0dmDLfkiT2QWXQJgQczEPAVEUWnZxs
AH1RV/jeU+nByyKtoKOPmjNII2jSI8AtK26EH77D9MR51Xz4hqQfMyaUEiq70UAdSUzHOL+jJOCR
czCpzZ31uzQY1FP/g4uZCVW1fd4OBUwKZZheEuN5pA/cNp8N8zMQWj8eSr3an7nATeYmd0JPahvn
GZDZ4gmGCJyLZ9NnP4x8qL8K0kTCMC5Xno4hC31Ta60R9mfCjNgJTzAkNSKS77vigFet0TZQ2934
BmYo2X4VFMRNdbkk6Kqk8u3tDblsV97K33+AC/VNdmH05t6krZftVz94CulhwtgX51vt72bomah2
cQAEDS2t8vCB8Bbr6iZI0LxzsP2VifKonpTxvIwV/G5uFTEO+azW20muGD/tDwvJ98/oxpnfvH+8
8ovZpfl2i94189uuOHYHGgPSmUsb4i7OEnV2wSekoPUokRqahE3axQE/WeUSXHTa5O2417n6KcKD
rPfvgryepjS8N9Wm4AiItlmULJtillGQIJDYl1bBauBeGf+BLXd779qVKfRhyZCeJ6tLKRcXDmmt
a18+7yIE365TXQYo4HTa7Laf3kyDUs/H2ThyMpS7OJgag4CgxsJHZsKRMqzqqTnbSMzVFEwif9mm
DOufExn5Fls1m3QTgUVRX5t9WSffLXzExIOvg6JStt6B1RsaZABCU9QoPTL7pqfpinCMfLAGDD/e
VQepnx9fwhxRf88W7VoVudE7MbUWRmWpi6q+lEZdEHuIo/UYjIDAB2bnoSMVDdUPjHgz6/XvY+jf
jgUdwrCPyQN8o5no8w1OGY4ELfKLyWI+iQ+BNtkwhaJ1lOkhxsBSPWDdaZKwdID9jIQ5qOigvusW
P2udR8JMi6m8qjm2wLF7ePUh5jj+qxXIqAD/xUzpSQS6VF7xZIkp4jGyF6FwQd9M7sGUTpSP9teI
OU2oa3UWNbgRlxXXP6eBu3jMauWzVtWsdoxJYV5vfaX/U59VWznfka2Yc58pMl/8j0I+PUy4c9fk
VNIXOLKduVSGvx1OC3Yr5Z6LdYjcR8hlry6hCtdcE9d2jrXivXoyhhyfIIHLCCrlgm0fNxTUh0c1
MrHwniHMxd86q163ryTa71ZKh5M34bD7tVcVivTVwwLcAYvW2ldJZIL5DCQHhoFXG7o84AZWqey1
SPMQ1CLnnoO3/7fIsh2aipT9YyA9iwqxJyFWo3Q8jDtsGfshQE9NczbKXdw82jRZvkxeBWVHCYOU
OcbFzYPI/+Xt9hrn5fvrSXOk5j/knSu9POc8MOZxUO9409OiDbGhjC7D+bTy+eVl6nc7qtWVnPmE
e+336EjQo8snR4l46wqJa4EwtTplMADwGu6Qgxa7Pkz8+ooOiwMhSPrxA2glvZAs7LYjz7okaNpJ
iUG3/dbDqr56eIwE0VyncwRGEdVna+ubEvnrfZVfzYui2vAAj0P7F7aTfL4yrhpIDrdH0ps1bTL0
AUBdMjHwS2AAHRH53fzgHb+7yBShqAcftCaKtYF5dV/SU08REqbkHS35HbPo+qum7b5UgxEkba4j
hB4mdbr/HDPPKpm9B7JWrYneyX9PRWC7APVZC52xP8JsIYhULTSR6Q2iGMkhiTGZFDrEW41V0bvo
g9C/KCnkVuaxWC6Wd/XaXbygFoZqVQfOrEiGSdSC/tUD997Yj0qRj3orSGl0tqfdTlgvKqhy6fyt
cNKl8l4Mv4XC7nZ9imx2j8RyrcUwZdJMAXqdVeTAX9QNzqe9nHJvd1I4EHWpPYCQOPlEhPMuBPUS
JuRpmTm1IPtD5VVIqZk1XtHXZcH7onFrXC4qibYBqr+H3FO9FmrPm0eqV9cO8jZbPTji/ZaC8xez
x+BZJjAm25VH965HNIC4p+Pb5nO8AEvUdrUu6xJ3P+OtiY1BeLMjr8MT9KIwH0NiDylpOtKxfb+C
vF+3lzjL2zKloWo80ZX8Y+ZRRcKpaMkbpMNcxUM0DmSla+W/PRijOxKv642d+nwrRu1uqbIkIXh1
IuInYRoSuJbfBri14rGrjGW4gjQeCWSJfW212yG5slAGMabW2TpWbokE3IQ4MWI8/eG9YGq4DLV0
TI/eIcCdyxLeEflFm34uywFpjiZEzeutcbwZvgb/MXHFl91vynHnQGCkTuRqKRxccCH0npbCg7jg
epxG3pPN7CLM+s+Ty7VRyjdwdm37+jcRy9z2HY2nKwve6v9S1Y7Awqucw2n7LkfhCwp7aEtBcVVL
Uuae1TI6kDBIljtYse/emwpXOWY2FWxxssbLKTFOjaEUzZmmlDgTD1dhpCvPVJjjprImSj3DE20F
4nJ0svtvzHII7zP+EgAhPgH11IxApaVAhgCIoXIjEV3suu+a+1PAgz1ExVs1rXb5l55zVtKJg+zV
Nk2MYv2/+viF291inytq00vbsVrW1fsWtCdfODkUR7MAsVQKlIXjnqNQBrKhEf7CQbVY0kWDTL7/
T2vBRgraBTG7/9uSu1XObF9GfZAhI9m/G0i/WllQoQLmz6eZMbrXtjCtGvCxfC1liKR7jUn0poXo
C+S8s0BlIwwtjInUYUGKfGRUAE0kQt8xhX0IzHFkUHvhurPHW+wOQnMGmkRF7wzmQds41sTabrnK
+2+uskZb/YR3qE5QPSWt1VSbKNGHjR5A3Nk/LamYJPMuBrOC2CF7iGUNSZVdgrQpBXezvmh50jm7
PkJXfpXojVn4IyeHsQq33A44DrebADhcTI1CIyB/KjcwEcEOiKyfVzs8+UCp+IeRhUuOv9e+OwG8
C9guJ1g2XYyYcR7W32fsn4XfjqXr2HIQVxqxANFB4HukRrSLUIo1/RXy+7K7M6WFzMnqYAUIVLiI
0jlarcDhjCagaBZknzzzP+hmL84/6pcUf+dctifTdhj5INmxdDGm9cT/RiRhJRG+JgZ10taRHh+q
3Z+mn9u1V1gSRlCLM+H4hBONsDFhxaKK6jG9ggjcRNc+N7V66paPv0o1ZOXSsKQ3kog4c36fl3d4
drEP4HY+fSaag8XGM4AXcwhtZqlhsnXSUooKJniivWtw8jFoQ4WMklyzgeAQA9Oj4UW4UDhG9c1c
gJZNIPb9Q9SSNsmHHwPAFMms5JIzlkR5FxUWliy6KwxaG4qNT9VF6hrkOZZqIup9QIgMHUv06Xdz
dr12LboQpctDEbYvtbMSfVUn5qm+4JpNpSomVHBQRs5JhDjWkSPXx/zalAgWkwNfgZ+psf8VcG2H
B773Tm2nsoFnOxPCmxRG9KhoGNEk9FwavDPSGkqhzXF3hJXYOpwaQKKOJaGHThkCr8lhXvpcScjJ
TLMEz4B1ohZc7DlGmznjRRvZLg2Mp24Q2R4K+XwcF7uBSlZN9xk4uapu0EATthJz7t7hsPllqA9n
W1++AroVmkrCFYL/wvBPsaI/mFVqZJKuaRatyWbpnNmveWEq3k6dvOH9E2AI+LItp4rJaA7kDUtF
/XUJep+7UHTwh001JosSKjsWF/GbDfziIIR5UnuSdOuyHNgKCdQgHcPhtVHjrP17Zi70RkAUcg3d
49nuVwBWKrtFQxM7VBjGgCnbkPsUyhzT3ICm0Vlrn6xK/MhDo7S6EW2ujQgy25wRwaYcvcapWC1J
M92+YpKkK6LrNVajMdcEbMeexxjzJE/lJPVeWI/eDykSiwnLarLae4ZepOr5Xv3MwsXVEtnk9IR5
w8ftub8HTo8FBCAZn7W6QXtcbe0ZIio/gy3kQeEnhhC8h5NCVuSmdE+Qy4gbWnSqQvY6xsFybK2Q
Y7e9iMiA5B82v2C4QHh6crGcTUYojrQ/OryCEIAJK31a3wYxFbjyEspGmIKhjJMtDYHNIUF2qQeD
FYnvdyWTlXEQAFFLLCsFpf+fp9TTz2Is5CYrIk28RGkLLnnV0RI8HCTZ47KSagDCFm1+gCiS7+jj
4yd5h/MiOVtQE2abvnfSZVgRiuMUTTNflfD1jMzDHGG6Pus/1n26U59KRKtKXh2nMzQIpPWL4bxN
Hxj/gt9bevYVS6mGQcKx84Ch1zFCopXW2dsAxBbBYL2jUaFjQD6WCQo9EZCaQZSX7gI/HHWYbauR
Gi9ydOrQby3NJzumAuBgpwzLlq4xXXr63VbYjWcDzcTXC98eEqQ7FdnL5OOy3/JKCP8fDjed+OhR
xvKTdnaJOW4EhZI0oEPvcqYIbR5qI7N2bSzgf3ZtR9ubHNctI08nlDSWIwZUHMbek5XGYY7xrGcJ
HyOHCk5EvQakUT4+jkIjii+goKn+6bG/JUzYYrGMKTI9NXXdpsTpd+uLauECA6zkM8fk5ix9Rga6
LP6yvKO6jw99veXu/dcK8N2u4qTnlqLlZIAi/oUTnmg+A5U9eizvOesyUANuEAu5SdfOvqCMoxr6
HgGp9qWQKtD86mHd5klnHy7D0RB3mV2WG3kTJKgelYa3blkHnrXeaBneMpWrnOMK9Az+R9mpsHsX
YyYz5wUmoejsoZHutFLbmtS0xKhWRyeZ8PsfxlJsx0DrvSpWCTn64AR4OgV2jpI9SRJOB+0l/xzi
NWbOUbgCMzngJa5QdRHGQznAyOjpEnytsiHeAjtwt4oVz4vRA/xDTf1CJaocOT2evnMXBNXsWxvY
Knc5TMTnFfKurXt+e09CrO24mID6BJrHIxGZxWnI0v3ILoxmY/wCrg/DPoGkJYEYd8VHuy1fKYN7
MxE6/z5yonLI6RbVfo6pMYiAYaj3xElhxOoro2U+v1JRNCzekr2tFvJRhnN0/xMyehNJatxQzOrL
XTRva5gE7bYCLokwCElljuNlLEEFcqIiQVxTxlkomXxxzngsv6PtALur4C+K+R2DPcM91E+AOjAC
o6/xEF5kui1PWp+ZNu+SsyANF8E1aYo/6pTjSWfDZFH1PjmGbbBVtglzkvR6YsZ6gEv/CaAwU6pQ
Z4OBFBDWcQ++b1PnmjJIU4vAHwIlARW1wow5idgz1MI8jsWxCXypwWNj9qwPQEAkN63yBapPsRAn
e4ViuxU/xVQplVl209WtXJF+XjXxaHktfL57KPAyo/xHVEh4o3sDK+JPzD7rMa+9PIY4X8m34hMV
L1bShb+LENR05gJlJVRaxggsVGMoYpnqChVTLtOr8cUxjIMpwP+qqqFGW59ekMdT/RxCyot661pM
Vg69WAFCOrAkibvF5JUrw55Ja2tBsL2REXiaswEZ97ZgV9HfqS8sLdk4huEU8pVz4uB4lRY/vpdf
lS1MYvDAF8XMSEI5pBtlTjksAO+BPosLfrikmPFYTtg0mF5HODV+cCpNeUpaPDMNiNiIy5EO1ehh
ZMYwvsYZEoiLdt+U+SwzZMLog5ONJ9NiHCh6Oq0iQ6wOHFmcarpgFkP3jsM4dUkrY1j+s7Qh9vZJ
CmtJp6yB6YAvp/BETmuoVD14GpVxgmobijdYoW3OIXv6Hb/tfnf9HmdFJMBh+7jWqDmmt2Ydmtd8
a/37xa7CHQEgD5Is/IQQcR8cEnqePC9bMnfWW7cl0wH6UYGxW/nPu185G4ugKTWvT/cv7jAeHYc4
fdfhCz9blMz9tWkwe4aPbGH92RkZRTZUIcS/NvKJAcoOX1klB5NaP4xK9w5PidMd5CgSbfQBrWkl
2G2bzldxnHugWRQ6CyN6HbYtMuh3LuvfBRMjcf9b6Muon0yGCTUhVALGbb+LFsDySm4Hq/gT0M5K
IOhOz+HATN16RfAqGv0/4c7DHlHB/Gjs1oFRI7T8YWXxktOl+prWE+HSrw+3PK0J2j0dTVoryi3P
MtDDi+0Yby8TYJsmW9lClKAgaNYs/nmS2pekSg2kp90ev7oq7W9Cz/hyp+KG80ctHoAAYShLDfOi
38PLu6jxrwPkEaKKQXqjaFxr9jsnsgOlXP8lj9Fudz6cJyz6d86BmXx6g+Kq0N7PfhTBkcC8I5Dh
b0j/5uQeSX31BA0F1aSMLVwjrZbRUBFGs1FD+7b+OShTNfjp1l2exP8oVrkZ98OHhawLizLibINA
qtihzFwD3L9gDgz+UPohiuB0N1/Sd3ZmxD+AyVQqO6TFgwJwxSuQrkFIrTbr4/lpH40EeB53jrwi
a1twno3FVvZqHphMWEoniR6QSZn6FuV8UnwzhfbBjPHLRzad7F7iw4bt6zwH72ZLaSwXX55jLEbd
aSHIljaFl4p8/lCeT36uYLRs5H8rrKvr+QsdkJZH0RwSdaVqCEiyBxlBXjLIdt1OU+s7JLvTvq/E
1O19ADx1DEuZjSkVmiJZoemQSVQ335yF6CSpy4tUvslnxJp61PacaFZ8olTz0RLymhEhCbbiHWmY
9t49ugSlZKD+URY8poAEBFId1pOwXhjn2XXhmrGb6RJ45sUI+aLBu7ZMj0S3jw9AKJDWCvWeg3kV
i0vCbEOXQT4YqDJtfNb/C9VwZVVvOuY8JgE6VWDx3BGEIc0us0tLDgG00mmFblJPoZHaWeOSep+B
HINIdy/YvAhJh/4TYaSIWt4Fyx5SJf3Heqk/nCDJSFrCgGjXsKvYnwRczTdl5yGkMA1twSoJvlWq
oARvqMcESgVj/LeJb9e+vkAMTAHTNqpHU+DPpsMkz+rjvX9S4AaVzDaCprN6iv5+e/WWQqJ9p9CC
79urcJvotaz/UsnljSraR5GYIUad5tYv/2YK4HdRU50FWtVjIM6jpL4ga4DWhryciYgiuVxpuxRg
5tXo2GqP062UTnxvsWpl7+0H8jdkRWFfKI8JZNpxJOA98a/xXe4RriRvKqPfTeRx7MejtKsdcRNq
AzCDdbE2ZwzMbsNq9bQFmmP8NIZZ8Ydkyv1hu6A5a5GaP1BSMr3H7yQXrI5hM7Kd8WnEjs+c+G1B
o5nqOvznfaB2wZmsEjIXaJAdCJPXX7HjWYW0IVseUtyWrfBljPbwM10tpuAxVPvwBl9ijd/mzswz
idxEUb4q6DkZm7QlbdLe/pQ5HdwUJc/wlMCdS2Ybgwn7SBFB6KaRAMvzzcZdKhctylm8hXBWCdsa
O/erS6FUt6efCWyu2nNA1aSoPlojK11GkhR8rcmaKblv0XEaWLjVUonJgpjvRuB+kznjVcbCOHY5
/n8a+chZZZICbsgFEC5hpnYfXh/8wv/zKo07vmIAi1aObiNE5HkdDwThh+oFiGnmVCxV7x0HGRo8
DUwv5PgrAOKiRoWnAArCiF/n4v1mOOwT9PvB4s5Jt1AGTn/e9/HxeJftQFwmZrWoDeqHp14Kv7jy
IrBZxBzKmQMLX0Uuzg+sBqZwohi8s9aVxbIfDDG5Ea0mlY2rHOaDYVM3KacbUeY4oNXwYaUUNi07
r1MYxDy3tciOqmp0HoZPjyHwuQaMOUtptNFr1ajHDv4I8gjn4kRF5qCuMoTb9pg6hGG5s8eJFSAL
7HpKvugisBPihnbQvVvS1WhGKxQQRQ8otTWdSeFk/PXI8b+LKxut/XVU81ziGJyhcfqsWTo+/VGY
s67xoY6yUhOBxwxKLrZzQCI7yvXMUn1yyTF0txsSxiIViisY2AwpO3heAVXPQYDJa69fIY1A9s+A
mU+eHj1wWn6AD23x31OXSOO3/3kor4sAXfE43x5GXLgRXhCStj5oO3viHibEOJwqr+fXSpsMQe9p
WDuX4i4l0ibVvfKS6RlXqk7Gta4PnWox5z6i/HraT/ijB95tv0ejnEqvNUzSZvSQYI2rokjzmz70
PAm7uD9W6q/SCtMQWZuS2K1PlpMXBuA/wxuldLanDNr2YZUhm9M8SaR6f+F+HN2xrJ9+Y4DWNp4j
Y0Z3yzEDUU51GixM6vBg9+8qmOfHaPjC9vH94GBEWVuulEwGhPMdLW3s+fLt2ySE7oRyukEBSYXT
HPYXnYlOGoe2ug1U8EpcRxCGj+qPB5N6BSrTgM6zZrcHaLFaZuJuaS7/y2HNaX3Ob+f+NWcUjqtE
LrfI+0+40x7B0dC5cFpuCLDtpC73FDKBAljc2COV+H/3Cq2p2Mg2Xm8K3YFa9M55DT3NpOpxt3gp
3lmJWs0lv6nIPousL4kVIYxRvXT819/eqweOC/9pufEzxMHDJ+CD19hrfUqPYNR0aecifgJBQ1Ya
B1ykA8XF0/x7Grls6lF8Tkc4C8xzkdiIYFN9xeGE7eJW/RSaU3OcszN+2XCN0ZOdJldMCHtwOv8G
6wbh/oa1+eOp0CBkOCs/2klrcDw8VPEd58psxqrefyE3dPT5ucDCbLEvioTgQvshXrxX3t+D4+93
JcViOBm7ZllnVWkw91QX7O1/NDP7aqpaqfvde1sQ+lojdaDWoTEVXvh+BD3pr1HGUBtS5n8ofKb0
cOZw8Ocsvx6XVuQ5rZ2AhJResPtTW1tb64pwDG3Ks7IC9JKiMp4iMczVARm+s00h9NUC0eNJBGzy
zIN2JyyiWuu3TNd9wV8OMdeuVapW0QAwYSGLOhruiFsmw8H2fg+QgpX3zIaBn6Js+xZ1OGi0lC70
494iUnfhsERDEoqrDkHDg8QqOS523HSjg6HZdF0SuI7Fs8FOwen6xLcLRAq5t4ZHG8gfltyCNg6V
XOs30PHU4tU31ns7aV3S3BBpAmS6Z7wGXG7pyzjbet2TelqOAH2WyFui46ofTSl2akASqZiN5u5o
hhj8eAHG8R+DBhdy2Orwpo0U0Phe08KlUzzsdyr2Q3soeHYodI+2R09xrpIi/dzsMiUMMjClkUnM
ckQZGvHZKGUrBOhSIc5aDi2MEP6Owoq8iQPi6vH5lH/RZmfm2li66g+DkcV9iLv14IFCP1Mzs1t0
0+JwVGpruaLQ5LAxCInVcu55ui64tFy0ErJYcxYR5MCKJl4JLrUFDlFlMjVfb9lxUfmn22mJ4toB
bDqAGRbPhIcSpxKXuv3U3vjzpm2wjRz8rn97r4h28fMG1TyA2voFkIZ+7XEu1HjnZTedMiBOyTuP
RoPBjK23kfqeCMogN4EC0DYADIig5X7SZE5WZ2wyMlRUaB17dH1Hqb1EkR68wlsFiqUiYbaVSMus
/ATtEosBM2DQzVLSXlW+aOkZ1pfWo9F13s5252L/3y2AE1kQ6J7Q4ycAxkkEF581su4falkOIfYj
dSwA8KjnqaDaA+zJ0TNTf16JLbAg4K290E6PWudy0Hs1NDGfpIHaWUkmcMaxiVD/oVQWsJae1J7n
wsS62o5Q+nUlnnxMjygWoUGPkDXmwsbFzBdDEznC5A07n1CZTPbVx+vnPLflV9lqXsh8fuq+jION
wxfxp8y+St8YmaCZzhAhVXbB+x951rRkhCT0NTJkuN48Ix3tL6Nx6BccIoNOrtd7C1gImYZvJ5rW
nD+hlOOzdf4onkHsZxt8FqxU1cqBNTcbFryceHDH2XZBIjTBcnXdTZGEytr19oe6UdNhCZzzkP6v
pAn1Dd+GwdPHGGNaMrs6hfeB1VYKPOZTITNfVR/CV3rgtJYq9BdrwybSlm8ejF05eZGizUYSLbOX
HMCc5EdAmAGosGz/vFjifM/7fbMsrdtEphalwX0d5EUtNarct2gK3Kgdp8Otl7XQ2u0DpovK9ZLp
VMOBX1rZrpPt93ASxRVSXByKRXBJyAIVBcD78jgwgZF8HCaLM7zSj27nBdQZQKFYXgo+88FrQnTW
ivDPZCbjIP/vZnlhJTDE5LDGYtK0U6TYN+apJsHSzILv5L1z0Zr1v5LGHPAtKlLTAm8ojzzsJDeT
t5oUq90gRaFKHDGTeBRV3I7+MEZtRI16aiaosEOc9satWgOqfcuyZeuLVtquC/byOVOLe7nk3Idi
L6p990OGjNI8D4X+JRc/2LtGHtAm7WjAMI1A1w/uhjH+fJm00yl3ahW4GRnXeJTH5sAyCCwHn16/
8gWZdxXDjSjnkw6p/SO33Vt82Nr3IHrQ9fVfPN0BCiMaKYRnTTHlPZVVY6xAct7zRWksvzUy+y29
MIilMfbQHV7fNAWT/9K6D+U7e7OydBqdTb0o6DeHRT+0S5flTQKNQkJbDSlFmxfMnD1LKtHW1w8x
yznmAaclCeymQ0lAf9HntvPKfZuzn1j446r8HlRfl27fFleA1SAk4STM4e7c36XBmv7KYj24vzd4
3xIU1KUV/fpMtZlBVTI5z6hTICurwa7C2Qu+k3hhjqg2/vaacP4xofshks9Vs0Z2nG4c4fZOBrH6
1YO9G6MjoWpwCmWy2oyAtdZYdV1fSsBPD+tE1n4+B+ZLZqhWlGbVRlhDKPJCaj8smLRa5FvgvbQz
5rA0hfNCH/mzrNSNYFzg4Ayj6HBvYf41hC3gT4uNePscJfNDgmOzlwLu6wF25TKiAeHObo0IuH3L
vqOwlPO8kPLtBSnp5OT6ynsbXQP1T7NUMhIkhkx9aj8XMgnAaNNz8Ms6WUmOIdc+3RfUH9r0r1PT
kEQwVjfx/ORz8SeHF9qB8ZPrilyGKSee3tLRZjmqWw3tzce+lrr6KNQG0Qpk0XoGkFcWnHbuEH0Q
xyGtG+rvqdsiMMhOkedHwiGofIxIK//+xOJe4YGLDH1z3h5I2BDn2Nz9ItV2ou7+pM0lCOsIFdfl
oUiq6JdGpOym3zjz/ktGMY1gztyEXwws+/LjDxtiK2pDIjhflSC1jY34k+S3M2y2y/Wl25P4RFAv
DbuPldp0uvHlT94jqr6LUJ0OSneoJ5MgStsXFwVzkrNdlnB7bL9asScuVPaudfXvO3VIHokBTvyH
2YV9rw4fWDxEqQRm0HG0l3SMCBkeQIsPnXamcTKg0r+xvtmIFEshEeGa2pEG3rmWGM+CUAM2ExNK
Am4bvdArpssxsIjeo+WFFUWprHUAH/Pbn7zCrRsFtFfqteA+ewdj95ptXV6qSY2H5Rnukls1LeoK
+opcg609zraOqZXxPV1Vp/H1NQuwstWOjK0t8tQGfPBfOw69IHzsh4PtPDrEQMnCzDBkDq2z9zJr
RwkI/KCDy5sCQNIpBINFCSG5iIhfAIKq3nxuxhHr2ypbJ37u8jZqJq4qT9+Eifn2DK10gjqm6GWz
og/zNhxXZBgrYiEwOmRGPQiu7s+FFN7Y+VeDaADj4drnQfgljn0Ufemc2WSPBtB0z+loUUAiMB02
whRGIu4S+GIwuGGa+n5NPCj47qo9KgE3b7Pvlq+QSI3CgBAwn4Mp9Uu+xcDpODSQhiePq7+PqcWi
zhCgv6KxwZ7OKZpOxPUc1axvmUN9soZspv99ptwmnOZ0tk/TScqPY43bmqOThzB/C53qh1EXMSI/
9CINDthx4L7tJTezCxEsL3sjNdsB+XKvemsWzons/I/xu3oqldGE8+gwrPKShipKpkDzWNrPjTQH
nqvasKBpjLiX+Jihk/RK6zZn/UoECl1ZH8c8egzrlaRJi7a7mJtHkXSW2C1kSHVFMHtl6tqCdLQK
B4oNcY5ZVgqyhweXGzoeZ6IMONWBwagbYowzV8MrnAa56fvuw9xp5cCQOBBPJmnLI9KNjlE4XaHy
/d6+mZj2wi87X1WwLl631YoOI19I++N+uAkzsWW8WAkXgkdWPiKVZxUNpu9nco+CCnovadwP2KpA
2vj44VG1jeJzyQ2IzJ8lQjU3+1psztRHPnPGfDTVZi+44HrFRUdngqbD0fiT0lEC3FpFmcjBtS1o
Q6oSCr1rGlV0tCr1hywh5hmu0nZrGDJjr0oKLq/V4dEd1j8Au5IW3dcGoDtUx/RB487W6k9O49Kx
iyZLhqBd6zk4BdnTDDhNE8baPSsk+gfXJGJKypobetbf9ih7X8+i+0dS+c4zNfyit51jrIkZf66n
eg==
`protect end_protected
